// X0Y1, W_IO
`define Tile_X0Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000100000110000000000000000000000000000000001110000000000000000000000
// X1Y1, LUT4AB
`define Tile_X1Y1_Emulate_Bitstream 640'b0000001110100000000000110000000000111001100000101001010011010000000100010100000001100001000000000010110000110000110100000010000000010100000000110010000010100000000110010000010100000000100011100001000100100000110000000000010100001100110000000001000000110000110000111001000110000000001000011011010000010000100100010011000010000000100000001000011111000001111000001000000101100001000010000001000000000001100100010000000000000100110001010000000010000000100000000000010100000000000000010000000010001100011100000011010101000011000000100100100000010000000000001110011000100100000100000000100000000001011001000010000000000000010100000000000001000000
// X2Y1, LUT4AB
`define Tile_X2Y1_Emulate_Bitstream 640'b0000000000000000000000000000100000000100010001000000000000101000000100110001010110000100000000000111100110000111001000100000010000110001100000000000100000001000000000000000100110001100000111101001100000100000110101000010100110001000000000000001000001010010110000100001000110000000011001011000000000110000100000000000000000000000000000000000001100101001001001001000000101100000000000000010000000000000000000010000001000000000000000000101000000000000000000100000000010000010000000010000000000010000000001000011100100000011000010010111100010010000000000001000000101000001001100000000000000011010000001000000000000000000000000000000000011000000
// X3Y1, RegFile
`define Tile_X3Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000011000000100000010000000001100000001000000111000001010000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000100000000000000000000000000100000000000000000100100000000010000000000010001100000011000100000110000000000100011001110100000000100001010100000000000000000010000000000000010011000000000000000000000000000000
// X4Y1, LUT4AB
`define Tile_X4Y1_Emulate_Bitstream 640'b0000000000000000111001000000000000100000111001110001010011010000000001000000000000000011101010100111110001001001110100001000000000100001100001100100000100110001010000000000100110100000100011100001100000000000010100001110011100001000000000000101010001010101110000010001000011000000100000011010000000011100110100011101000101000100000000100010000000000000111011100000000100000000100000001111000000000001000000000001000000000000000001000000111010000001100000100000001001100000000000010000000000100010010011001010000100000000111000010000010111000000000000001010011011100000000000000000000110000001000000010000100000000000000000010000000100000001
// X5Y1, LUT4AB
`define Tile_X5Y1_Emulate_Bitstream 640'b0000000000000000011010110000000000100000101000000000000000011000000100100001100000100000000000000010000110000000101000000011000000100000000000000110100000101010000010000010001001001000100100000000000000101000100100000000010110000000000010111001011000000100001000011001111000001001011101000000000000100010000001001100001101000000001000000010001100110000100100001010000000000000000001000000000100010001000100100000011101001000000000101000000110000000000000000100000001100000000100011100010011000010101111000000000100001000100011000111110000000010000000000110001010000111001000000000001001001000000111000010000000000000100000000000100001000000
// X6Y1, LUT4AB
`define Tile_X6Y1_Emulate_Bitstream 640'b0000000000000000111110000010000000000110011000110001100001000000000000110101010000000011110110000100110000000000000100001000000001010101000001110000000000000001010110000011100000101100000001000000001110101000010100001100011001010000000010100001000001000011011000000001101101000000001101111000000000000110011000001111110100000000001000001001101000011100001010000000000011000000000011100001000000010101010011110000000011010000000001001100000101001000100000010011000000000000000000011100000001000110000000000011000100000101000000110100001000100000000000111011011101000000100100000000000101110001010000100000000000000000000000100001100011000000
// X7Y1, DSP_top
`define Tile_X7Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001001001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000010110000110011101011000000000000000010011011000000000000101000010000000000000000000000000000001100000000110000000000
// X8Y1, LUT4AB
`define Tile_X8Y1_Emulate_Bitstream 640'b0000000000000000000010000000000000011011101001110000000000000000000000110001010000000001111110000000000110000000110000000000000000001100000000100000100001000000000010000101010100001101001000001000110000000000010100000101100110000000000010000000000110000001110000010001101101000001000000011010000000000110000000010000111100010000000010000000001100111100001000000010000001001101000001100000010100000110110000011001010110000000000001110000000000000000000100000001010000110000000100001000000001000000111100000010000000000000011011010101100000000000000001001111000111111011000100000000001001110110000000000000010000000000000000000000001000001001
// X9Y1, LUT4AB
`define Tile_X9Y1_Emulate_Bitstream 640'b0000000000000000110000001000000000100000001000010001000000000000001100100000100000100100000000100000100000000000000000000011000000000000000001100110000000000110000000000111000000101101000010001000111000001000010100001111011011010000000000000000100001010001001000010000100101000000010000100000000000000100010000101000000011000100001100111110001111010000010010000000000000000101100001101110000110000101000000000000000100000000001000000000000100000100000000000000000000010000000100000100100000010000011100001100100000000010000111000111000000000000000000000011001001101010001000000011001110000110001001101010000000000000000000000000001100100000
// X10Y1, RAM_IO
`define Tile_X10Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y2, W_IO
`define Tile_X0Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000110000000010110000000000000000000000000000000000000000000000000000000000010
// X1Y2, LUT4AB
`define Tile_X1Y2_Emulate_Bitstream 640'b0000000000000110001001000100000000010001000001111011001010000000000000000100000000010010000000000001110000110000001100011110010000110101000000110100000010001100010100111010011010101000001110001001100100110110000010100010100111011000000100100000110000100010000000001100000000000001000001001011000001000000000100000000000000001000010001100010001111000000001000100000000011001000000000100000000000001101100000111000010100111100000000000100001110000000010000000000000000100000011000000000000000000000000101011001010000000000010101110011100100000000000000001001000110010011000000000000000011000001000111111000110000000001100100001110010000100000
// X2Y2, LUT4AB
`define Tile_X2Y2_Emulate_Bitstream 640'b0000001000000000010001100000000000001010101000100100100000111000000100000000010100010010011100000000010010000001000100000110000000011100100000101100000101000100000110001010000000101101000000001001000100010010010100000001000010001110000000000100000000010100111000010000100010000110000101100010000001000001011100010011100011001000001000000100001100110100110000000000001010110011000001101000000100011010011010000000000000000000001000010111111000000000100000100000010000000000000100000010110001001100001011001000100100000001100100100011100110010010000000000100000101010001000100000000001100100000000101110000000000000000011000010111000100000000
// X3Y2, RegFile
`define Tile_X3Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000100000000000000000000000001000100010010000000000000000000000001111110100000001111000011000111100100010000000010000011111101010110001001111001000000000000011100110000000000010110000000000000000000000000100000010000000000000000000001000000000001101000010000000100010100000000011000011111010010000010100000000010001000000000000000000001110000010101110000000000000000000010011111100000000
// X4Y2, LUT4AB
`define Tile_X4Y2_Emulate_Bitstream 640'b0000000000000011100100010010110000000001100000010000001010010000001001101000100101100001001000000100000010011100000001010110000001100100000001010001010001000010001000100110000011100000111100100001000100000110010001001110000101010110000000000100000101010110111000001000000010000001111101000011000000010001000000001100001001110000001010001000001000111001000001001000000100000111100001000000110010000010110100011000111110000100001000001011000001000000000000100000001101010000001000001000110000011110111100010000100000000010000011010001101010000010000000000000100011100011000000000000001010011000000110110000100000000001100000001000001000110000
// X5Y2, LUT4AB
`define Tile_X5Y2_Emulate_Bitstream 640'b0000000000000000001010001100000000001010000001011011000000000000000100000101000001101111111110000101010000000101101100000000010000101000100001000111110000000011010000000000001001100000010000100001000000100111000100101001001100001110000000000000000010010000110000010001001110010101110000000000000000000010010100111100001100101000000000111000011011000000000011001000000100100000000000000000100000010011011000100000110010001000000001011000001100000000000000000001010001100000000100001000000000000001100000000000100000000011000110000010000000000000000000011000001100000100001000000000000010000001100100010000010000000000000000000000000100000000
// X6Y2, LUT4AB
`define Tile_X6Y2_Emulate_Bitstream 640'b0000000000000000101000001100000000011110101001011001010000111000000000110000100100110000000000000011000000001100001001110000000001101001100000011001100000000000011000000000000100100000011000000000000000000101000000100110101101010100000000010000100000010011001000000001011010000010000011001000000000001110111000001010100000000000000000101000011101000000001010000000000100010101000000000110010000000000000010101000000000101010000000000000000000000000000000010000000000000000000000010000000001001000100010000010100100000010000010011110000000110000000000011101101010001110001000000000000000000010101110100000000000000000000000000000001000000000
// X7Y2, DSP_bot
`define Tile_X7Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000101001110000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000110000001100000000000000111000000000000000011000000000000000000000000000000
// X8Y2, LUT4AB
`define Tile_X8Y2_Emulate_Bitstream 640'b0000000000100000100000000000000000011110000001110011101001111000000100000000110101100111000010000001000000001110000000001110000000010100100001001001100010001000000110000000001010001100010011000001010110000111100101101100010000001100000000000100000000100011110000000000010110000000010000011000000000000111110000000100001010011000000110000000001110110000011000001000000100100000101000000111010000000100101000110110001010000100000000110101000100000000100000000000000000000000000000011000000001000000000000001000010100000001000110000010000000000000100000011110001001011000000000000000001001010100011001100000000000000000000100010000000100000000
// X9Y2, LUT4AB
`define Tile_X9Y2_Emulate_Bitstream 640'b0000000000000000000000100000000000100000101000001001000000101000000100100000000011110010000010000000000010000000000100001011000000100000100000110010000000000011000000000100000010101101000000001000110000001000000010001101000011010000000000000000101011010010000000000001100001000010000111000011001100000001010100000011100100101000000110001000001111000000000100100000000001001001100000000000100000010001101000001000000001010000000000011000000000000000000000000000000000100000001000000000000000010100000000000011100000000001000101000111100110010000000000010110000100101011001100000000001100000100011000000000000000000000000000100000001001000000
// X10Y2, RAM_IO
`define Tile_X10Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000
// X0Y3, W_IO
`define Tile_X0Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000000000000000000000000000000000000000010000000000000100110000000000000001000000000000000000000000000000000000110000000
// X1Y3, LUT4AB
`define Tile_X1Y3_Emulate_Bitstream 640'b0000001100000000001000000000000000011110000000000011111000000000000000000000100010000011111000000101000000000010100000000010000001100000100000100010010000000110010000100101100000001000011100000000101000001111010000010000010000000000000010000100010000000000110000000000101000000100000011100000000000010011001101001100011000000100000100000000001111100101000001001000000011011010001100001000010100010110011000101000001100000100000010010000110010000000000000100000000000000000000100010100000001011001110011000000100100000000100001010011000000000000000110000000001000000110001000000010100010111100010111000000000000000000111000001000000010001000
// X2Y3, LUT4AB
`define Tile_X2Y3_Emulate_Bitstream 640'b0000001000000100100000100000000000000100000001010101111001000000000001100011000110101001000000100000000000001001000100001110000001000001000011100111100100010011010100000010110000100000110010000001100010100001010100001000010000001100000000100000000010100000000000010000100010001001100001000000000000110100111101011011100010101000000100001000010100110000010000000000000001000001000000100111110000010101010100010000001000001000000000000101000000000000100000000000000110110000100000000000010000000010010100001011010001000000000001011111000000000000100000011000011001010100000000000000000001101100000011000000000000000000011000010000001010110000
// X3Y3, RegFile
`define Tile_X3Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000110101000000000001100001000100100011000010000000000000000000000000000011111011011000110000000000000000000000011101110101100010010011001101000000000000000011000000000011001100000000001011010100000000000000100001100000000000000000010000000000001101010001011100110100001011101100000100100001010000110000000000000000000000010010000001010100010000000000000000100000000000110000000000000000110000001000
// X4Y3, LUT4AB
`define Tile_X4Y3_Emulate_Bitstream 640'b0000000000000000110100001011000000011011110001110110111011100000000100001000110100100111000000000011010010000010011000101110000001101001100001100010100000010000000000000000101100000000110110100001001000100000000101001110000100001000000100000000010001000100001000001000010010000000001101010000000000100000010101101111100011001000000000000000010101100001010011001000000000100110000000100110010000000001001001001000001000001100000000101000001000010101000000000000001101000000101001000000000000100100011100000000000100000000000000000100001100000010100000000111001011000101000000000000010000110010010000010000000000000000000001001001100000000010
// X5Y3, LUT4AB
`define Tile_X5Y3_Emulate_Bitstream 640'b0000000000000100011111100001010000010010110000000110100000111000000001000001000000011100011100000001000010100000010100001000000000001100100001111100010101010001011000101000000000100000100110100001100000110001000100000100011100000010000100010000000010000000000000100001011000010000101001100000010000100110011001011111001010100000000000111001010000110101010101000000000100110000000000000110110100010100001101010001101101000000000000001000000110100000000000100000001101010000000000000000000001001101100000000011010000000001000000010000100011000000000000010010101010101000001000000000000011001010101101000010010000000001100000000010100011001000
// X6Y3, LUT4AB
`define Tile_X6Y3_Emulate_Bitstream 640'b0000000000011100100000000100110000100000011000000110111010000000001100100000000000011100000000000010010001001000100101111000000000000000000000000110000100100010001010100000000101100000100011000000000100000000000010000111010000000000000010000100011010000000000000000000100000101000001000000000001100001001010100110111000010110000001010111000011100011100010111000000000000100011000001101000110000010001100010000000000111101000000010000000000100000000100000000000001000000010010000010100000000000100000000001000000101000011000110010100000000000010000000000101100001001000001000000000001100010011100000111000000000000000000000000000000101100010
// X7Y3, DSP_top
`define Tile_X7Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100001010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000100000000000000001010000000000000101000000000101100001011000000000000000000000000101000000000000111000000000000000000000000000000000000000000000000000000
// X8Y3, LUT4AB
`define Tile_X8Y3_Emulate_Bitstream 640'b0000000000000000001011101100000000000010010000100001000001110000001100001011100001011100000110000100010011001000010100001110000001100001000100000000110000000101010000010110010010001000000000000000000010000001110000000011000000000100000010100100100001001001110000000001101100100000000000100001000000001001001000111100001000000000001100000000001101001101100101000000000101010000000000001000000000010101000100000000100101000000000011000000000000000001000000000000000000100000000100010000000000001000001000000011010100000001110000010101010000000000000000010001001000111010001000000000001010000100100000000001000000000000000000001100110010000000
// X9Y3, LUT4AB
`define Tile_X9Y3_Emulate_Bitstream 640'b0000000000000000000110001100000000000000000000010000000000000000000000000000000000100100000000000000000000000000001000000011000000110000000000000000000000000000000000001000000000001100000000000000000000000000110110000000000000000000000000011100100000100000000000000000011100000000000000000000000000001111000000000000000000000000000000000000000000010001000000001000000011000000000000000100000100000101000000001000000000000000000010000000000010000000000000000001000000000000000000000100000000000010100000000000010000000000010000000101000000000000000000001000000000110000000000000000001100010000000010000000000000000000000000010110001000000000
// X10Y3, RAM_IO
`define Tile_X10Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y4, W_IO
`define Tile_X0Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000001000000000000000000000000000001000000000000000000000000000000000
// X1Y4, LUT4AB
`define Tile_X1Y4_Emulate_Bitstream 640'b0000000000011000000001000000000000001011111000101000000000001000001000011101100100110011000110000001000011000110100000000000010001101000100111000000100000010011010000000010100100100000000111000000100000100110010101101100000000000000000000100100000001101001000000011000000000001001101000011001000000000001001000011000000000101100000000001000000010000000001010100000000011010110000000000110110000001000011000000000001000101000000000010100000010000001010000000000010000000000011100000000000001111010000101010010010001000010110100100000100100000000100010001100100100000101000000000001000001000011101100000000010000000000010000010000000110010001
// X2Y4, LUT4AB
`define Tile_X2Y4_Emulate_Bitstream 640'b0000000000000001010000101000000000011000000000010001000001110000001000001100100000100000000100100110010100100000000100000110010000101000100010100101110000010000010000100100100010100000110000000000001000100000000100000100001001010000000010000000000010001000110000011000101100110000000000000010000000010010010010010000001010000010000100000000010011000100010110000000000010000000000000000111010000000100000000011000000101000001000010001001100000000001100000100001001000010000000000000010000000100100000010000010100001000000010010000010100010000000000000011000011101011010001000000000000001001101101000001010010000000000100000000000001000000001
// X3Y4, RegFile
`define Tile_X3Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000010000010000010110000000000000000000000000000000010100101000100000000000000000000101001000000110001011001001000111100011011001100000011000000100000100000000011000000000011110011000000000000000000000110000000000000001100100011001011000010111111000000000001101110000110001001001101110000001001010111000000000001011000100111000100000000000011000000000000000001110000000011
// X4Y4, LUT4AB
`define Tile_X4Y4_Emulate_Bitstream 640'b0000000000000100011100001100100000011110000000110101110001100000000100000000010011110111000000000011010011000001110100000110000000101001100001100111010100001000000100000010100100100100001100000000110000100010110100010000010010000000000000001100101111001011000000000000000110011000000000000000000000000000010101011000010100000000001100000000000010010000000010000000000000100111101111000000010100000000001100000001000000000000000001110001000110001000000000100001000110000000000000000000000000011000000100001000000001000000000100101100010100010010000000010110010100101000101100000000000010000110110011111010000000000000000000101000111100000000
// X5Y4, LUT4AB
`define Tile_X5Y4_Emulate_Bitstream 640'b0000000000000101110001010000100000010111110000000000000010001000000000000000000000001100011000000000000000000000011100001000000000111000000011000010010001011101010000000110110110000000010100101000000100100000100101011001000010000110000000100100000101100000000000010000010100011111100011110010000000000111001000001111011010000100100000011000011100110000110000100000011000010111000001001001000000000101001000010100101100000000000001100101011110000000100000000000000100100000000100010000010001001110110100001000100000000011100111000111100010000010000000010011100010000100001100000000000001001000000101000010000000000000100000001000100100010011
// X6Y4, LUT4AB
`define Tile_X6Y4_Emulate_Bitstream 640'b0000000000000000001000110100000000000000001001110011100000111000000001101011000111110010111000100110000101001100001000011100000000001101000001100000000000010000001010000100100010100001111110100000100000000001010001001101010010000000000000000100000011000100111000000000000001001001101001000011000000010001000000000000000111101000000010001000001111001001010001001000000110001000000000000001100000001010111000010000100000000000000000000100011011001000100000000000101000000000000000000000000000001010001010000000010000000000001010100000000000000010000000001011101001001000000100000000001010000010010001111010110000000000000000000001000000000000
// X7Y4, DSP_bot
`define Tile_X7Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000001000110000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000011000000000111000000000000001000000000000000000001000000000000000000000000000000000000001000000000000100000000010000000000000000000000000000000000110000000000
// X8Y4, LUT4AB
`define Tile_X8Y4_Emulate_Bitstream 640'b0000000000000010000111000111000000000001010000010100001011111000000000000000000110000101001010000100010000001110010101110110000001011001000000000001100001000011010110000100100010000001000000000001110100000000000010000010000000001101000000000000111000010100001001010000011001000000010100100001000010000010001101000100011001101000000101101000000000110000000010001000000000101110000001000101110000000110010000100000001110001100000011010000000101000000100000000001000000000000001000001000000001000000011010110000000001000000000010010111000010010010000000011010100011000100000100000000001001001101001111101000110000000000000000000000011100100000
// X9Y4, LUT4AB
`define Tile_X9Y4_Emulate_Bitstream 640'b0000000000100001100000000000010000000110000000010001110001100000000000000011000000000001110110000001010000000000000000000000010000000000100001000010000001000110010110000000000010101100010000000001001110000000000101011100010000001001000000010101000001011001000010000000111000100010010011110010100010011111000101000000100100001100001000111010000000010000100000001001000000100001001101001000000100000111001000010000000000000100100011010100000000000000000000000001000001000000000000010000000000100010110110000011000100000000110100000100010000000000000000000000000101100100100000000000100100000000011101000000010000000001100000000000011010000000
// X10Y4, RAM_IO
`define Tile_X10Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000010110000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000
// X0Y5, W_IO
`define Tile_X0Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000010100000000000000000011000000000000000000000000000000000000000001
// X1Y5, LUT4AB
`define Tile_X1Y5_Emulate_Bitstream 640'b0000001100011101000000110000010000000000101000000000110001111000001101100000000011100010001000000001110110000101111001011100000001101000100000100100000101001000010000000110010101100001101101100001100100000000100000010111001110001000000000100101110010010000000000000000011100001000110101111010000010000101011011000000011110000000000000010000000111100000001101000000000010010110000000000110000111000000011000010000001011001001100010000110100000000000001000000000000100000000000000011100000000011000001011000000100100001001000010111000000000010000000000000111011001001100001000000001000000111100010000110000010000000000110000001000000110000011
// X2Y5, LUT4AB
`define Tile_X2Y5_Emulate_Bitstream 640'b0000000000100101110000000000100000010101010001111001100001000000001100001000010000011001111100000000010010000111111000110100000000010000000000001001000000000010000100100100001101000000000000000001110010000110000100001000000100001101000010000000000000000010000000000000101110000000010001000000000000010001100100101111111100001000000101011010001000100100000000001000000001000001000000000110000000001000000010000000101010000100100001100001000010000000000000100000001010100000000000011000000000000100000000111101000100000011000110001000101000010000000000010100001100000010000100000000000010101100000001100000000000000000100000010101010000010000
// X3Y5, RegFile
`define Tile_X3Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000010000010100100000100000000000000000000111100000101110000000001000000000000000010101010100010000000000000000000000110010100001101011000101001100000000100000000100101011000010001001000100001000000000101011001100000000000000000000000000000000000000011100101011111010110000010000101111000000000000101011000011000000000111000000110001111000000000011101110111000100000000000000000000001100000000000000000000
// X4Y5, LUT4AB
`define Tile_X4Y5_Emulate_Bitstream 640'b0000000000001000100000010011000000000110000001110011101001111000000000000011000001110011010000000001010000000010101100001110000000110000000011000111110001000011001100100010101000001000100100000000000100100000010110000000011000000100000010010000110000000110001000011000111001001111000110000011000000000111010011000011010001000010001010000000000000001001000011001000000011001110000111000001010000001111100000000000000000000100001011110000000000001000100000000000000000000000000000000000000001010000001100001000100000000010011100000100000010000010000000011100001110100001001000000000000011101010100001101000100000000000000000010000000000111000
// X5Y5, LUT4AB
`define Tile_X5Y5_Emulate_Bitstream 640'b0000000000000110100100010000100000000000001001110011100001110000000001100000010000001110100110000111000001011000000000101110010000001000100110010001110100100011000100000110100000100100110000000001010000000001100000001101000000001110000000011001000100100100001000000000010010101000100000010000000000000001101101001111100001101100001001011000001100110000110010101000000001110001100000001111111010010100001111000000001100000100001010110000000001100000000000000000100111000000000000000000100000011001111100001000100100000010001010001111100000010010000000010010010010110000001000000000000010001000010001100000100000000000000000110100100000010000
// X6Y5, LUT4AB
`define Tile_X6Y5_Emulate_Bitstream 640'b0000000000000001000100010000000000010111110000100001000000000000000000001000000000010000111000100010000011000000000001110000000000000101000001100001100001110000001010000000101000000001110001001000000000100111000000101011000110000000110000100000100001010000110000000000010001001000000000011000000000001010010010011011110000000000000000000000000000101000101010001010000010100100000000101111010000001000011100111000001110010000000010010111111100000000100000000000110000000000001000011000010001011001110010001000010100000000001111010100000100000010000000011001001010000010000000000000000100001010110011000000000000000000000000100000101110000000
// X7Y5, DSP_top
`define Tile_X7Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010100000000000000000000000000000101010100000000000000000000010000000001101000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001011000000000000000010101010101010100000111100000000111000000000000000000000000010111001000000000000110000001010000100001110101111000000000000000000000000000000
// X8Y5, LUT4AB
`define Tile_X8Y5_Emulate_Bitstream 640'b0000000000000001000000011000000000001111111000110000000010001000000000000000000001101001000000000101000000000000000001000010000000000001100000000101010000010110001000000000000011100001010000001000000010000110000001001001101010000110000000100001100101010000000000000001000011101010000001110010000000010001100010000011110000100000000100101000010001111001110001000000000101101101100001001000100000000101000000000000101100010010000000111000000101000100000000100000001000000011000001000000000000000100001000001001100001000000000000000000100010000010100000000001100001111001000000000000000000000000000011010000000000000000100001001000000100100010
// X9Y5, LUT4AB
`define Tile_X9Y5_Emulate_Bitstream 640'b0000000100000000101001010000000000000000101000010000111010000000000000000000000110101100000000000000010000000110011000001000000000000100000111011100000000111000000100110000001000100100100110001000000000000010110000001111111011010000000010011100000101000011001000000000010001100010000011010010000000001110010111000000001111010001000010000000000000010100110110000100000000101000100000001001010000010100110000010000010101001001000011101000000001100000101000000000001000100001000000000000000000000000000000000000100000000001010000000000100000010010000010010001011000111010001000000000000000001011000001010010000000000000000000001000101100000000
// X10Y5, RAM_IO
`define Tile_X10Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000100000000000000000000000111100000000000000000000000000101100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000
// X0Y6, W_IO
`define Tile_X0Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000001000111111100000000100100010000000000000000001011000000000000000000000000000000000000
// X1Y6, LUT4AB
`define Tile_X1Y6_Emulate_Bitstream 640'b0000001000000110100001010100100000111110000000110000110000000000001100000000000000001000110110000010000001000000000001011000000000101100000000000111010000010000000010000110001000000000010010000000100100001101000000000000100100000010000010100000000000000111110000100000101100000000000000000000010000000001001000000011000100001100001000000000000011100000000000100000000011010011001000000001000110000000001111000000011000000100000101010100010000000000000000000000010100100010001000000100000010001100011001000000000000000101000000000010100000010010000001000110000110011011000100001010000000111000100110000000000000000000111000011100000000100000
// X2Y6, LUT4AB
`define Tile_X2Y6_Emulate_Bitstream 640'b0000000000000000000100110000000000001000100000100000010000100000000100000100110110111100010010000001000011000110001000001000000000001001000101010000010100001011000001011010010001001000000000100000000010000011010000000000010100000011000000101001010001000000000000010000010111000000000100100000000010001010001100100000000000011001001000000010000000001000000011001101011111000000000000100000100111100100000101111100110110011110110100001000011100000000001010011000010100100000101000001100010000000100000010100001000001000001000100000010111000000010000000000000011100011001110000000001000000000000001000000001000000000000000000010000000101000000
// X3Y6, RegFile
`define Tile_X3Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001001100010100000100100001110000101000001101111001000000000000100000000000000111100010110100001100111011000000011100010001000110110001111111100100011001100001000000000000000001001100100000000000000001011000000000000000000000000100000000110000100100000101101001000000101110000000001001001010000000000000011000001000101000000011111000100000101000100010010000100000000000011000000001100010000000000000011
// X4Y6, LUT4AB
`define Tile_X4Y6_Emulate_Bitstream 640'b0000000001000110111100001000100000001011111001110011101001010000000101100101000001110001000000100010000110000010101000000010000000000000000000100110100000100010000000000110011000100001110000101001000000000010010101000111010110001100000010100101010000110100000000000101100010000000010001010000000001001100000100011000001000000100011000000000011011010100100000000000000000100010101000001011000000110000000010100001000010000000000001011000111110000000000010000000111000100000001100001000000010010000000011010111000100000000000001000000010000010000010000001010000010000000000000000000001110111001010111110010100000000000000000001100101101101000
// X5Y6, LUT4AB
`define Tile_X5Y6_Emulate_Bitstream 640'b0000000000000001000000100000000000000001000000100101000000000000001101101000010000001100010010000010000111010100010000010110000000010100100100010001100001101010000010000010100110000100001110001000110100000111000001000100001011010100000000000000000101010010110000000000001000011101110011010000000000000010000000110011010000001000000100100000000111010000000010100000000010001000000001000001000000010101001101110000010100000100000010110110101100000000100000100001001010111000100000010000000000011000000000001010100100000000000101100100100010000000000000010001001111001110001000000000001100000100100001100010100000000000000000000110001101011000
// X6Y6, LUT4AB
`define Tile_X6Y6_Emulate_Bitstream 640'b0000000000000000010110111110100000000010111001000001000000000000000000001110010111111101010000000001000010110000000100111010000000011100100011100110000100100011000010000100010001101000110001000000000100000011000100100100000100000110000000111100110010010000110000000001100101001101101001111011000000000110101000011110000000000000001010000010000110111001111001000000000001011000000001001001100100000000100110110000001100001000000010110000000100000000100000000000000000100000000100000100000000011000000111001011000100000011000001101100000010000000000000011111011010000100001000000000000101001000010001000010000000000000000000110001001001000000
// X7Y6, DSP_bot
`define Tile_X7Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000110011000000000000000000000000000000000100000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000110000000000000000000000000000000000000000000000000011000000000010000000000000000001010000011100100000000000000000000001100111010000000000001000000000000000000000000000110000000010000000000000000000110000000000
// X8Y6, LUT4AB
`define Tile_X8Y6_Emulate_Bitstream 640'b0000000000000011011110011000010000000010000001110111111010000000000000001001110000010101011000000111000111001001001000100000000001100100100111100010100101001000000100110100110001101100010000000001010100000000100100000100000000001100110000001000010001100000110000010000010000100000000110100001000000001000000100101101011110001000000101000001100000110100010001001000000010000100000001000100010000001000000100100100001000001100000000010000010100000100000000100000000000000000000001000000100000010011010000110001100001000001000000101100000000000010000000011010001111100000010100000000001000010110110000001001100000000000100000101001001110101000
// X9Y6, LUT4AB
`define Tile_X9Y6_Emulate_Bitstream 640'b0000000000010001001000010000000000010111101000010001011011011000000000000101100000100111000110100001000000100000000001001110010000010001100000000001000000000000010000000110100110000000001000100001100110000000000100001001111100001100000010101001000101000000000000000000100001000000010001011000000000010001000100010000100010010000000111100010000011101000001010001000000011001100000000100101010000001100100110011000000110001001000010001001000000000001101010000101100000010000000000011110000000000010100001001000000100000000110100000001110000010000000000000110001001000011000100000000001000110100011011100010100000000001000000001111001000100000
// X10Y6, RAM_IO
`define Tile_X10Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000000000000000010000000000000001000000000000000000000000000100000000000000000000000000000000000000000001000000000001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100110000000000000
// X0Y7, W_IO
`define Tile_X0Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000100001100000000000000000000001000000000000000000000000000000000
// X1Y7, LUT4AB
`define Tile_X1Y7_Emulate_Bitstream 640'b0000001000000001100011111000000000000110011000000000000000101000000001110000000010000001000000000010100010010010000000000000000001000001000000110100100001100100000000100110001010001100110001000000000000001010000100000000000000000000000010010000000000000000000000101000101011000000011001010000000000110100000101011010001010010100001010000000011100000000110000000000000010000110000001001110010001000110101000101000011110000000000000100000100000000101000000100000000000101000000000011000000001000000001010010010100100000000000010001111000000000000100111010101001110101000001000000011010000000000000001100011000000000000011001010110000110100000
// X2Y7, LUT4AB
`define Tile_X2Y7_Emulate_Bitstream 640'b0000000000000000000000000100000000000100000001000010011010111000000101000010000110001100100100000110010100000010001100100000000000100101100000001000110000000010000010110000000100101101110001100000101100000000000101000100001000000100000100001000010000100001111000001001000110100000010010011000010000100011100000001011011001000100000000000000000001000000001000110000000101000000001110000110001000000000001110010110100000011001000001000001011100001000001000001001101010110000001000000001011001100100010100010011110010011000001110100000100100000000000000001001000000001111001000000000001000000010001000000000000000000000000000111110000101110000
// X3Y7, RegFile
`define Tile_X3Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000100010100000100100000000000000000000000000001000000000000000000000000000000000000110111000000000000000000000101000000010110000000011001110101111100011110011000011110000000000100001000100001000000001000000000000000000000001000000001100110010000000100101111100100010001101100010100100100000110111100101000001000001000001101010000100000000000101000111001000000000000000000000000000000000000000001000
// X4Y7, LUT4AB
`define Tile_X4Y7_Emulate_Bitstream 640'b0000000000000101000000000100100000001000101001111110010000100000000100100000010001100101010010100110000110000010100000000010000001100000000000000000000000010000011000010010001000000001000000001000000100001010000000000001010010000110000010000000000000010110111000011001101100000011001000000000000000011111001000001100010111100000000000001000001011010101010101000000000101011101000001000001100010010001000000100000000101000000001001110000100010000100000000100001101110100000000000000000011001111000100100000000100001000001110000000000000000000010000000000111100000000000001000000000001110011000001101001000000000000000000000001100110000001010
// X5Y7, LUT4AB
`define Tile_X5Y7_Emulate_Bitstream 640'b0000000000001000100111000000000000000010001000100000000010101000000000100001010001000111000010000101110110000001000100010110000000000101100000100000010000001000011010000101111000100000000101101001010010000001000100000001000111011100001000010000100000000010110000000000001101111010000011010011000000010101000100000000000000100000000111100000000011001100000011001000000101000011100000100001100000000110100001001000100010101100000001111101000110100000010000100001101100000000000000011000000000010010000010001000100001000000000110010000101010010010000000011011000100000111001100000000001001001110101001000000010000000000000000001000101100100001
// X6Y7, LUT4AB
`define Tile_X6Y7_Emulate_Bitstream 640'b0000000000111000111100110000000000000010000000000110110011111000001100001000110111000001000000000101000010001111000000000000010001000001100000100000000101001001010010000100110011101100010001100001101000100000110010100111001100001000000000010100010001001001001000000000001101000001001010100010000000000001001000101111100100011000000100000010001000001100000101000000000001010000101100000011000100001101010010010000000101010000000010000010000000110000100000000000100110110011000000000100001001000100001000001000100000000000010010000000000001100000000000010111110100000000001000000000100010000100010100100010100000000000000100001000010000001000
// X7Y7, DSP_top
`define Tile_X7Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110010000000000000000000000000000010000110000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000001011000000000000000010100000000000000000101111010000000000000000111100000000000000000000101000001101000000000000101011000000000000000000110000000000
// X8Y7, LUT4AB
`define Tile_X8Y7_Emulate_Bitstream 640'b0000000000000100000000001100010000001000000001010000000000101000001101100111000010000000000010000010010110110000001000000000000000101000000000010010100000100010000100010010000001100001001010101001100100000010000100101011000110001000110010000000001011000001000000011000001100000000010001000011000000000011000100111000011000011000000010000010010001001001000010001000000000100010100000000110000000000010100100000001010110000100000010010000100000010001010000000001010001000000010000001000000001100010101100000001000001000000010011000000000000000000000000011101000100000001000100000000000001010000000111111000110000000000000000000000001000000011
// X9Y7, LUT4AB
`define Tile_X9Y7_Emulate_Bitstream 640'b0000000000000000110000010100000000010001000000000110000010000000000000000000010000000000000000000100000101110111110001100000000001110001000110001001100000100010010110000000111001100001100000101001000000000000010000001101000101011110000000000100001001010010110000000000100000110100110001000000000000001001001110001011001000000001000001100000000010000000100010000100000011010100100000001110000010001100001110001000001010000000000011010000000110000000000000000010000000000000001110010000100000101000011100011011000100000101000101010100000100010010000000101100000100000010000000000000000100001010100011000000100000000001100000101001001000000000
// X10Y7, RAM_IO
`define Tile_X10Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000001000000011000000000000000000001010000000000000000000110000000000000000000010100000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000010000000000000010101100000000
// X0Y8, W_IO
`define Tile_X0Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111100000000000000000000000000000000000000001001000000000000000000000000000000000000000000001000000000000000000000000000000000
// X1Y8, LUT4AB
`define Tile_X1Y8_Emulate_Bitstream 640'b0000001000000100100000000000000000110101010001010000000000000000001100001000000000101010111000000001110010000000111100001000000001000001100000000100010001000111000000000010100100100000001001000000000000100000000000000000011000000000000010000000000100100001001000100100100100000000001100010000000001110100010000010001000101100000010000101000011111010000000100100000000011000000000001000000100000001100011010000000000001000001000001001000100000000100000000000000001000011000000000010000000000000000010100001001000100000101000101100011000000010000100100001100011111110000000000001100001100000010100001010010000000000000010001010010000001000000
// X2Y8, LUT4AB
`define Tile_X2Y8_Emulate_Bitstream 640'b0000000000000000000000010000000000100010010000000100110001100000000101100000000001010111010010100000010000001001010100100000000001001000100001101011100100100011010010100000001000000001111000100000100000000100000010000010101000000000000000100101100110110100000000110000000010010000000000011000011000101001101010000000000010110100001000001010100000011000101000000000000010000001000011101110100010000010000000011110000110000000000011110000110100000001000000100010000110100000000000001000000000010000001110001110110001000010000100001000100010010000000000010001010100100000011000000000000001010000011000000000000000000000000000010000000011110000
// X3Y8, RegFile
`define Tile_X3Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000110110110000000000000000000000000000110010010000101100000000000000000000000011001110011000000101000000011000110001111011110101111111111000000000000000000000110000110000000000001001101000000100000000000000000000000000000000000000001100111000100000000001001100100010001101010000001001011110111111000011011101110000000000001101000010111001000000010000000000100000000000001100000001010000100011000011
// X4Y8, LUT4AB
`define Tile_X4Y8_Emulate_Bitstream 640'b0000000000011001101011000010000000000000001000100111011010111000001100001000110111010000000000000100000010001111000001110100000001101100000000001001100101100010000000100010001010000001100010001000011010000000110000000101000010000110000010001100010010000000110000000000000000000100010010100000000000000000001000101100001100000000000100000001000011110000110000000001100000010010001000001001000000000010001010000000001010000000110000011000000110000101100000100000000110000000001000001000010000011010000000011000000000001000000010000010110010010000000000001010000011011000000100000000000111001100111000110000000000000000100000010000010100010000
// X5Y8, LUT4AB
`define Tile_X5Y8_Emulate_Bitstream 640'b0000000000000000000110100000000000000000000001100010111011111000000001000011100001110001000000000000010110111000001000000010000000001100000000100100100000000010000010110010011011100001001100000000010000000110110100001101100000000110000000111101010001011001110000000001101010001110000001001000000000000010100000101011101010010100000110000001101101000100011100101000000000000000000001000000010000001101100000000000100101000000000011011000000100010001000000100010011010000000010100010000011001001000001000001000010000000000000110000010010000000000000000001010010100011001100000000000001100011101000001111000000000000000000000010000000100010000
// X6Y8, LUT4AB
`define Tile_X6Y8_Emulate_Bitstream 640'b0000000000000010011000000100000000000110000001000110000000000000001000001011010110000100000000100100000001000110111000010110000000010000000100000010000000110011010000000000001100000000100100000000111100000010100000000000001101000000000000011100110000001010000000000000010001000000000101000000000000001100000010000010000000111100000110100100001100000000100010000000000010001010000000101110110010010011111000000000100000000001000001100000000010010000100000000000111000000000110000000110100000100000000000000000100000000010110100011110000000000000000000001011001000000001001000000000000001000100010011100000000000000000000000000110001000010001
// X7Y8, DSP_bot
`define Tile_X7Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000110000000000000000000000001100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000111000000000000010100000000000000000001010100000000000000000000011100000111000000010000000000000000011101100111000000000011000011000000001100000000110000000000
// X8Y8, LUT4AB
`define Tile_X8Y8_Emulate_Bitstream 640'b0000000000000000110000111100010000011110000000000000000000000000000000000000000101101010000000000000010000000110110000011100010001000100000011001100010000010010000000000110001111100000010001000000110000000000010001000100001000000010111010100000000000101000000000000000000000000000000100000000000000000000000110001110000100000100000000011000011000101000000101000000000000101000100001100110000000011010010010001000011101000000000001000000010100110100000000000100000001100010011001011000010001011100000110011010100100000010000001000100000000000000000000000101101010011010001000000000000100011001000000111010000000000000100000100111010000010000
// X9Y8, LUT4AB
`define Tile_X9Y8_Emulate_Bitstream 640'b0000000111000000000001000000110000000110011000000110110001100000000001100001000000001100100100000100000000000110101000001000000000100000000000100000000100010000010100000000010100100100011000000000100000000000000000010101000000000000000000000000110001000100111000000001110010001100100010010000000100001000000000110011000011010000001000100000010011100001010011001000000010001100100000000000000000000010011000000000000000000000000000110000000110000001000001000010110000000000000000000000000000001100000000000010000000000000011110000001100000110010000000001000111000001000010000000000000000000000000110101010000000000000100000000000001000100000
// X10Y8, RAM_IO
`define Tile_X10Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001000000000000001000000000000000000000000000000000000000000101000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000
// X0Y9, W_IO
`define Tile_X0Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y9, LUT4AB
`define Tile_X1Y9_Emulate_Bitstream 640'b0000000000000000101001000000000000010101010001111111001001000000000000001010010000010000010000100010000001100100110000000000000001000101000110001000010000000100010010100100110100000000000110100001000010000001000101100001000101011100000010000000000010001010110000001100010000000000000001110000000100001110000000011111000000000000000000000000010000110100100000101000000000011110000001001000010000010100001101000000001000000110000011000011101100000000000001000000000100110000001100010000000001001000001011000000100100000100000001000010000100000000000000101100100111011010001000000100000101001010001111000000000000000000100000010001000100000000
// X2Y9, LUT4AB
`define Tile_X2Y9_Emulate_Bitstream 640'b0000000011000000000000010000100000000000000001000011111011111000000000100000000010101000001010000010010001000010001101011000010000000001000000011110000001000000000110000100101010100000011000000001000110100001110010000000101100001010000010001100010000000010000000001000000000011110000010011000000101000001010110000000000000011110010111000011000011100000001011011000000001000010100100000000010000010001100100000000011100001000000000001010001010000100000000000010000010110000001001000000001001100000000000000011100100000000000101000100100110010000000000001111011110000011001100000000000001011111100001000000000000000001100000011000000100001010
// X3Y9, RegFile
`define Tile_X3Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000100100000000110110110000000000000000000000000000100001000100110100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000001001100000100011000100010000000110001001000000000011000000000001000100001001101000000000000100011000001110000000100000011001000000000001100000000100000000011
// X4Y9, LUT4AB
`define Tile_X4Y9_Emulate_Bitstream 640'b0000000000000100011001001100000000100110000001010011101001010000001101100011010000001000000000000101110110000001000001111000000001000000100000100101110000001001001001001100011000000000011100001000110100000001010001000000100011010100000000010100100000000011000000001000010100001000000001101000000000010000000000011100110100100000000101100000000000010000001011000000000100100100000001000000100010000100010111010001010000100000000011001000010111000100000000101001000110100000000000010000000000000000010010011000000100000000000100000000100011000010000000011111101110101011000000000000000100000100110110111000000000000000000000001000000100000010
// X5Y9, LUT4AB
`define Tile_X5Y9_Emulate_Bitstream 640'b0000000000000000000100111000000000011100000001011011110001000000000001000110000001101001000000000100000000110001001001011110000000100001000000011001000000100011000000110100000000001100011000000000000010100000010000001001110001010010000010000000100100000011110000001000100000010000000001011001000000000000010010000000101110011000000101100001110011101100011000000000000011100010000001000001001011000110011101110000101000000000001000110010000010000001100000100000000000010000001000000100000000000000000000000001000001000001000110010101010100010010000000001110000100100000110100000000000000100001010000000001000000000000100000010000100110101000
// X6Y9, LUT4AB
`define Tile_X6Y9_Emulate_Bitstream 640'b0000000000000011000001100100000000011001100000100000110001100000000000000000000001011100100100000000010000001001111101111110000000111000000001100011000000100000011110000100000000100000101010000000010110100111110011001100100101010000000010101101101000000110000000001001100010000001000011001000000000010000100000001111000101000000001001000001100000100100101100001000000100000000000000001000000000010010010010101000001101001000001001111000010010000000100100100000111111100000000100010000000001100001111011010000000100000011001100000100000101100010000000000010000111100010000100000000000011010110111111010000000000000000100000100000000010000001
// X7Y9, DSP_top
`define Tile_X7Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000001010000000000000111110000000000000000000000000100000110000110000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000001000000000100000000000100000000000000000000000000000000000000000000000001011000000000000101000000000000000010000000100000000111100000000111011001001000000000000101111000000000000000000000000000000001100000000110000000001
// X8Y9, LUT4AB
`define Tile_X8Y9_Emulate_Bitstream 640'b0000001000000000000000011100010000000110011000000110000000000000001100000000010000000000000000000010000001000001000100110110000000001100000000000001100101000011000000010000000000101100000001000000001110000000100000001100001101010110000000001001110011011001001000000000000111001000000001011001000000000000101001011000010000100000001100000010010000000000011010000000000000010110000000000000110000000000010000101000010100000000000000001000000000010000000000100001000000110000010100000000010001100010011100000000100000000000010000000100100000000000000000011101000111000001011100000000001101001110111000000000000000000000100000001000001010010000
// X9Y9, LUT4AB
`define Tile_X9Y9_Emulate_Bitstream 640'b0000001000000000001100010100000000000010001000110001010010101000000000100001000000011100000000100010000100000000000000010000000001000101000000000010000010110000010010000010010010001100100100100001000100001000100000001000001100001100000010010000100000000000110000000000100000100000100000000011000000000010001100010011000000001100001001101000011011101000100000000000000000010001000000101011000000010011000000010000001110001000000000010100000010000000100000000001101000000000001000001000000000111100010001010011000000000010000010100100000000000000000000001011010010000100000000000000001000111011001001000010100000000000010000001110100001000000
// X10Y9, RAM_IO
`define Tile_X10Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000001100000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000
// X0Y10, W_IO
`define Tile_X0Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001010000000100010000000000000000000000000000000000000000000000000000000000000000000
// X1Y10, LUT4AB
`define Tile_X1Y10_Emulate_Bitstream 640'b0000001010000100000001010100000000000000000001110000001000000000000000100001110001101010001000000010010100001001011101011100000000001001000000001001010000100000001000000100010000100000101100100001100000000001010000001110100101011000000010010000000001010010000000000000000100100101100011001010010000100000010100000001110000100000000001100000000110000100001101000001100011000101000000001110100000011100000010000000000101000000010001001010011000000000000000000100001110100000000000000001100000000000000000001010100010000001000000010100100000000000000000011000000100000110000100001100000100000001000000001010100000000000100000011010000011100000
// X2Y10, LUT4AB
`define Tile_X2Y10_Emulate_Bitstream 640'b0000000000011000100111100000100000001010000000000000101001111000000000000101100111101100111110000000010000000001001100000000010001000100000000000110010101000010011010000000010010000000010100000000100100010000000000000100001100000000100100000000010001001001111000000001100011001001001010000011000100100100001000011100000001110100001010101000010011101001000011100000000010011101000000100010100011001000111001011000001010000000001100010100111000000001000000100000010010100000000000001000100001001000001100011000010001011010100100100000100100000010000101001100110110000011010000001010001110011001100001010011100000000000000000001001101101000000
// X3Y10, RegFile
`define Tile_X3Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001000110010000000010000000000000000000000101101001000100100100000000000000000000001110001110100000000000000000000110001101100110001101101101000000000000011001100011000001100000000010000000000011110110000110011000001000000100000000000000000001010010100110001010011110110000000110010001100101101110000000000101100000110000001000001100111000000000100001010000111010000111011110000000000110000000000001011
// X4Y10, LUT4AB
`define Tile_X4Y10_Emulate_Bitstream 640'b0000000000000000000001010000010000000000000000100110010011111000000001000010110100010001000100000001000000001100010000100110010000000000100011101001100110000000000100110100100101001101101100000001001100000101100100001100001000001100000000111000100101000001001000010000010001100000000000000001000000100000010100100000100101001000000000000000001100110001000011000001100000000110000001000001000000001001000110100000001000000000110000001000001010000000000000001100000101010000001000010000000000110101010111001000000101000000011101001111000000010000000000000001001100100100011100000000000000100000100110101011100000000000000000000001001011100000
// X5Y10, LUT4AB
`define Tile_X5Y10_Emulate_Bitstream 640'b0000000000000011011000010100000000101010000001011111001010011000000101110101000100110111000110100100110010000000001100100111010000100101100010100100100010110000001010000101111010000001100010001000100000000001010100001001011011010010000010000100000001010011111000000000000101001100100001000011000000001101010001000000000011100000000010111000000011110000010011000000000011000011000001001001100000011011101001011000111100000000000101010010101100000100100000100001010000100000001001000000000001001000011101001010100100000010000111100100100000010000000000001011011001000110001100000000001101010000101000010010000000000000000000000111001010010000
// X6Y10, LUT4AB
`define Tile_X6Y10_Emulate_Bitstream 640'b0000000000011110100101111100000000000100000000000100111000100000000100001000000011010100010010000000000010001010100000101000000000100000100100100010000101000100010111010100000010101001110011000000100011000000000001100100011000000000001010001000000000010011001000000001011100100100000000111000000000000010000000000100010011010000000000101001101111100100111011010000000011000001100110001001001000010101010000110010000000000000000010110000100000001000100000000000000000010000010000000100010000010000000000111000000100000000000100101100001010010000000000001000011000101000010100000000001000000000100000100001110000000000100000000000101001010000
// X7Y10, DSP_bot
`define Tile_X7Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000010000100000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000100101010000000000000000010000000001110000011000010000000000000000000000110000000000110000000010000000000000000000000000000000
// X8Y10, LUT4AB
`define Tile_X8Y10_Emulate_Bitstream 640'b0000000000000010110001000000000000000000100000010000000001010000001000010001000010100000000000000011100000000010000000001111000001000100000000010100000000101000010000000100001000000000101110101000000000100001000000001000000010000000100000010000000001100001000000000000011000010100000011000010000010011010001000001011100000000100000000000000010011000001100000100110000100010010010000001000000100000001000010010000000000000000000010111100111000100000000100000000001000100000000000010101000000001000000001001000010110000100000001110111100000000010000000100000001001101011001100000000000111001101011001000000000000000000000000000000001100000000
// X9Y10, LUT4AB
`define Tile_X9Y10_Emulate_Bitstream 640'b0000000000000000000000100000000000000110011000111001000000000000000100000000000000110000001110000000000000000100000001000000000000010100100000000000000001100010000010000001000001101100101000100001100100000101010000000000100100001000000000000001000000101100111000000000000101000000010010001011000000010001000101000000001001000000000011101000001111111000101010100000000001101010000001101010000000000000111000000000001010000100000000000000000000000000100000000001100000100000000100011000000001000001100000001000000100000000000110010100100010010010000000001010000100000001000100000000000100011001010001000000000000000000000000000000000000011000
// X10Y10, RAM_IO
`define Tile_X10Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001100000000000000000000000000001110111000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000
// X0Y11, W_IO
`define Tile_X0Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y11, LUT4AB
`define Tile_X1Y11_Emulate_Bitstream 640'b0000000000110010000000000000000000010111011000010001001011011000000100000000000110001100001100100100000010000110110101100000010000011000100000100010110001010100000100010100000110001100000100000000000010000000000100000000000000000001000010000000000001100001000000000000000000001000000000000000000010000001000001001100000000000000000000100000000011010100000110000000000001000010000011000001010010000100000000000000000101000000001011000100010100000000100000000100000001100000000000000000100001010000010010001010010000000011100010000001100010000000000000001010100001011010000000000100000000000000100010010000000000000001100000010000000100010000
// X2Y11, LUT4AB
`define Tile_X2Y11_Emulate_Bitstream 640'b0000000000000010000100000100000000000000001000110000000001100000001000101000000111110001111110000000010010001000110100000010010000011000000000100010100001011010000000000110000110000000100000000000000100100000110100000000000100000010000010001100000000000000000000101000000100000001010110100011010000101001001001101000000100010000010110010000101111100000000110100000000001010100000000000001000010010100100010000000001101000000001011000101011000000001100000000001000000100000001000000000000011100010100010001010000000001111000010001100100010010010000000100110100000100000000000000000000001001100000000000000000000000000100000001100011001011000
// X3Y11, RegFile
`define Tile_X3Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000100000000100111100000000000000000000000000000010001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010101000000000000000000000000000000000000000000000000100011001100011010000000010001000110000001010000000000000000000000000000000010000100000000000000000000000000000001100000000000000000000001100000000000000000000
// X4Y11, LUT4AB
`define Tile_X4Y11_Emulate_Bitstream 640'b0000000000000010010001110000000000010101010001100010000001111000001100100101000101010001000000000110000001001100011000000010000000000100000011111000100000000000000010000010010100100000001010100001111100001010100100010100010101011000000010010000110000001010110000000000001100110000000011000010000000001100000100001111100010000000000100000000000000100000010000000000000000101110000100000010000000010110001011110000101000000000000010110011001001000000000000000000010000000000001000000000110001001110001011001011000100000000000100000000000000010010000000001010001001000110000100000000000000111101110000100010000000000000000000011001001101010010
// X5Y11, LUT4AB
`define Tile_X5Y11_Emulate_Bitstream 640'b0000000000000010000000000100000000001010101000100100000000000000001000001000100111111111001000100100010001001110010000001110010000110000000100001101010101010010000100000100001010000000001100000001101000000000000000000011000000001000000000000000010100010000110000010001100001010100010010000000000000011100010110110000101000001000000000000000001000000000000000100000011110000010101100000111010100001110001001000000100110000000000011111000001000000000100000000000011010100000000010001100000001000001101110000000110000010101000000000001100000010010000001101010111010000101001100000000001100000000000110001000000000000000000000010000111100110000
// X6Y11, LUT4AB
`define Tile_X6Y11_Emulate_Bitstream 640'b0000000000000000000010011000000000000000000001001011000000010000000001100000000000100000000000000010100010010000000101000000000000111001000000110000000000010100001000000100000000001000001001000000000100000001110000000000101000000100000000011100000000001100001000011000011100010000000001100001000000011110010010010000100101100000000000011010000011010000100001001000000110000010000001001000100000000001001001101000110000000100000000001010100010000000100000000000000100100011001000010001000001100100011100000010100111000000000000001101000110000010000000000100101001001010001000000000001101010000000100010010010000000000100000100000110010000000
// X7Y11, DSP_top
`define Tile_X7Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101001010000000000000000000000000000010000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000101100000000000000000000000000000000000000001000000000011000000000110000000000000000000000000000000000000000000010100000101000000000000000000000101110101101101100000000000000000000000000000000000010010000111011010000000010101100000000000000000000000000110000000000
// X8Y11, LUT4AB
`define Tile_X8Y11_Emulate_Bitstream 640'b0000000000000000111000111100100000000000000001001000001001000000001000101000010000000010000000000000010101000001001000000000000001011101100100010000010010000000000000000100000000000001011011001000000110000101000001101011010010000100110000110000000001010101001000011000011001000000000011011011000000001110000000100011100111000000000111001000000000010000011001000101000010000000000001000001000010000000110000010001010000001100001010011001011000100000100000000000010000110000000000010000000000010000011110001000000101000000100001000010100110010010000000011100001001001010000100000000000000000111101110101010010000000000000000000000110101001001
// X9Y11, LUT4AB
`define Tile_X9Y11_Emulate_Bitstream 640'b0000000000000101101101100100000000000000101000111001000000000000000000100000100010100010001110000000000000000000000000000100000000001000100000011001010001011000000110000101001000100001000110001000100001100001000000001110000111010010001010000000001000111010000000011000001101000001000011000011000000000001011000001011000100000000000110100000000011000000000000000000000011011000100000000110000001010100101000001000110000000000001000000000100110000001000000000000000000000000001100000000100000001110010111011000110000000001000000000001000100010000000000011111010110001110001100000000000100000100000001000000100000000000000000010000101000100010
// X10Y11, RAM_IO
`define Tile_X10Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000011111111111111110000000000000000111111111111111100111111111111111010101000101010101010101111111111111111000000000000000000101010
// X0Y12, W_IO
`define Tile_X0Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000101000000000000000000
// X1Y12, LUT4AB
`define Tile_X1Y12_Emulate_Bitstream 640'b0000000000000011101000011000100000000010001000010001000000011000000000000101000010000010000000000010000101000010000000000111000000011000000100000100000000000100010110000111001000000000100010000001100000000111000000000000011000001010000010100001000000100000000001000001101101001000100000100011000000010001001111000001000110001100001011000000010000111100110110000000000100011000000001001000000010011000100011011000011101000000000010101110011000000000000001011000000100010000001000010001000000000100001111001011010110000001000100001100100000000000000000001111001110100010000000000000000000011000110001000000010000000000001000000011000010000000
// X2Y12, LUT4AB
`define Tile_X2Y12_Emulate_Bitstream 640'b0000000000000000100000001000000000000000000001100000010000000000000000000011010010001000000000000100000100000010111101111000000000101000000100000111110000000011010010000000000100000000101010000000010001000000000001000010101100000100001010000000101001010000110000001000000001100000000001001001000000001100000100000000010000110000000011111000000000100100001110000100000000001100100000000110110000010101111000000000001101010000000011010010000100000000000000011000010010100000001000000000011001110000000000010000100000000011000000000100100000010000000000010000000001010011001100000000000100000000000000010000100000000000100000011000111100000000
// X3Y12, RegFile
`define Tile_X3Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000001000000000000000000000000000000001010100001000000100000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000110000000000000000000000000000000000000111000001001000001000000110001000000011001000100011000000000000000000000000010100000001000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y12, LUT4AB
`define Tile_X4Y12_Emulate_Bitstream 640'b0000000000000000101001011000110000011000100001110110010011010000001100000100010111001100010110000011010001100011111101111000010000010101100011111000000101110010000000010000101011000000010110000000110000000000000001000000000000000000000010000000010000001000000000100001110011001001000011100011000000101000000001000000100100001000001110000000001000110101000101000000000000000000000001100000000000010000100000101000001101000000000001100000000100100000000000000010000000011000101010000100001000000000001100001000110001000100000100000010000100000000000000100101000011010000001000000000001001000100010000011010000000000000000000000001000110100010
// X5Y12, LUT4AB
`define Tile_X5Y12_Emulate_Bitstream 640'b0000000000000000000011000100100000000001111001010111010000100000001001000000000000011011010010000001010001010010100101011010000000100000000110000010010000000000010100100010101000101000001000000001100000100110010000010001000001011000000010100000101010000110001000011001100011001000101001010000000000000100100101000011111001001000001101000000001111000001010010000000000001000101000001000000000010010101000011111000000100011010001001110000000000000000000100111000000100010000001000000100010001100000001000000001100101000111011100000001000000000010000000000000000100000010001000000000000000000010100000000010010000000001100000001010000001101000
// X6Y12, LUT4AB
`define Tile_X6Y12_Emulate_Bitstream 640'b0000000000000000000010001000000000000100010000000000000001111000000000000000000101100101110100000001000000001101000000000000010000011000000000001100000100100000000110000000101001000000100100000001100110101000110110000011000100001000000010010000001000010000000000001000000000100001000000000010000000000100010101101000000110001000000000000001100000001100100011000000000000001010000000101011000000010011000001110000000010011000000000110001000100000000100000100000000100100000001100001010000000110000000000011000000000000100000000100101001100000010000000101110110110101001001100000000000001011000000000111010100000000000000000100010001010000000
// X7Y12, DSP_bot
`define Tile_X7Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001001010000000000000000000000000000010001110000000001000000000000000000000001100000000000000001000000000000000000000000000000000000
// X8Y12, LUT4AB
`define Tile_X8Y12_Emulate_Bitstream 640'b0000000000000000110000000110100000000110000000000110000000101000000001010000000000001011000110000001000000000110100001111000000000000101100000000000010110000000011010000010101100101100101010000000100100001000000100100101100000000001000010001101110000100000110000000000110001100000001000001010000010000011000000001110101000110100000010111000001111000001001001101000000010001111000000000000110000000011100011100000001000000000000011010000100100000000000000000001000010100000001000000000000000111110101001001000110001000000110011000111100100000000000000011101001010101000001000001100001001100101101010110000100000000000000000000001000000100011
// X9Y12, LUT4AB
`define Tile_X9Y12_Emulate_Bitstream 640'b0000001000000000000000100000000000000000000001111000010001100000000001010010000000101000010110100001010000000000001000100000010001100000100001100000110001110010011000000000000010101101001010001000111010000111000000001101110111010100000000000000001011110100001000000001010011000111000000001000000000000000101000100011000011100000000100000010001011101000011011000000000100011011000000100001100000000000001010010000101110010000000000000100000000000000100000100000000001111000000000001000000001001110010001011000010100000001000011110100100010000010000000001010001011100011000000000000000000011100000000100010000000000000001000011000000111000001
// X10Y12, RAM_IO
`define Tile_X10Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010001000000000000000000001111111100000000000000001000000001000000000000000000000000000000000000001100000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000010000000000000001111001111111111001000000000100010000000
// X0Y13, W_IO
`define Tile_X0Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000001010000000000000000000000000000000000000000000000000000000000
// X1Y13, LUT4AB
`define Tile_X1Y13_Emulate_Bitstream 640'b0000000000011001000000000011010000000000000000000001000000000000001000000000100000001100110110000000010000110110001101110000000000101000000010000010000000010000010110000000000001000000101100000001000000000000000010011100001100001000000010000000111111000000000000000001100001101001000100010000000000000001000101100011000100001000000000000000000011100000000111001000000000000111000000000101000000110001011000001000101001000100001000000000000100000000000000001000000001100000001100000000100001000110000010011000100000000010000101001000100100000000000100000010100111000110100000001100000001001000000011010000010000000000000000010010000000010011
// X2Y13, LUT4AB
`define Tile_X2Y13_Emulate_Bitstream 640'b0000000100000000001000010000010000100010001001000000111011111000000000001101010000001010000000000101010110110001001100111110010000100001100100010011100011010010010000000110100111100001001001101000000010000111000000000101001010000010000010111000000000000101111000000001100011001000001001011000000000000000100001110000000001000000000000101000100011101001001000000000000110000000000000000000010010010000000000001000001000000000000000110000000100001000000000011000010001100000001101010000100000100010000000011000100000000011100011010111100100010010000000001110001000010010001100000010000011101000111110000000000000000000000000011010000001000000
// X3Y13, RegFile
`define Tile_X3Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001100000000000000000000000000000001001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000010000000100000000001100000000001110000011100100000000001010000000000000111000000100111001100000000000000000000000000000000000000000000
// X4Y13, LUT4AB
`define Tile_X4Y13_Emulate_Bitstream 640'b0000000000000010000000001100000000011110111001000010000000010000001001101011010100011001001000100001000000110110110100010000010000001100000001001001000000110000011010100010001100000001100000000000100010000000100100001001001011010110000000101101000001000010110000000000010000011001000001000010000000001000011010010000110100000000001101000010010000101100000010001000000010010001100000101111000000000010001001010000001010000100000001010100000110000000100000000000010011000000001000001000000001001000000001010001000000000011010000000001101011000000000000010110000111100000000000000000001001110110000000100010100000000000000000001110000100100000
// X5Y13, LUT4AB
`define Tile_X5Y13_Emulate_Bitstream 640'b0000000000000010011110001000010000000110000000000000000000011000000000001011100110000000000000100001000100001110000001110000010000000001000111000100000100111011000000000000110110001000000110001000000000000000110000011000001110000000000000011001110111001010000000010000111101010000010010010001000000011110000010000000100000110000001001001000000011011000000000100000000001100000100101100011100001100110011100100000001010000000000010011111000010000000100000011000000000011100001000001001000001010100010101010000100010000010000010000001100010010000000000001010000011000010001000000000000101101000001010110010000000000000000000000010010101110000
// X6Y13, LUT4AB
`define Tile_X6Y13_Emulate_Bitstream 640'b0000000000000001001100001101000000000000000000000100001010000000001001001010000000000000001000000000000001001000000001100000000001111000000100000001110001011011010000000100000100000000100010000000000100000000100110100000001100000000000000110001000000000000000000000000000101000001010010000000000000010100001110001111111100110000000010011010000100000000010010000000000010010110100000000011110000000001110010010000110010011000000000011001000000000000100000000000000000000000001000001100000001000100001000000010000100000000000000000000000110010000000000000100000000000000000100000000000010000000000000001010000000000001100000000111010000000001
// X7Y13, DSP_top
`define Tile_X7Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000001000000000000000000000000000000000100010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000011000000110000000000000000000000110000001100000000000000000000000000110000000000000000000000000000001101000000000000000000000000000000000000
// X8Y13, LUT4AB
`define Tile_X8Y13_Emulate_Bitstream 640'b0000000000000000111000000001000000101000100000000001000000000000000000100001100000000011001110000110010001000000000100001001000000101000000000000110000001001011000000000101110000100001000111101001001100101010010100000000010110001010000010000000000000001100110000000000000001000000011010111000000000000101001100001111001010100000000000001000011101100000011000000000000001111101100100000110100000010101001111000000000010001000000000110000000110000000000000000000001100000000000000011000000000101110010000000000010100000011110110000000100000000000000000011111001010001001000000000000000110000001100101010010000000000000000000001000001100000000
// X9Y13, LUT4AB
`define Tile_X9Y13_Emulate_Bitstream 640'b0000000000000000000000110110000000110001000000000100000000000000000001000010010001000011100000000101010000001000000100001001000001110001000011100100000000001010000100000110110001101100001011000001000110001000000101000111100001011100000010000000000000010010110000000000100101001000001001101000000000000001010100010011000000011000001110111000010011010101001110000000000001001101000001000111010000000001100000010000100101000000000001111101000100000100100000000001010000100011001000000000000011010000000100011000000000001001000010011100100000000010000000011100000010010010000000000010000101011100000000001000000000000000000000000000001001110000
// X10Y13, RAM_IO
`define Tile_X10Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010000000000000000000001000
// X0Y14, W_IO
`define Tile_X0Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000001
// X1Y14, LUT4AB
`define Tile_X1Y14_Emulate_Bitstream 640'b0000001011000000000001001011010000000000000001111000101001101000001100001100010010100000111110000001010011110100000000100000000000100001100001111010100001000100010000000100111011100100101100000000001100000000000010010100000100000100000000000000001110100000000000100100000101110111101110100000010000000000010010010101000100000000000000001000010110101001100111001000000000000010000000101110000000000000011010000000101011010100000000001000000000000000010000000100000000010000001000011000000001000110101000000000100100000000000100010110100000010010000000011110101110001010000100000000001000101001101000100010110000000001000000000000001001101001
// X2Y14, LUT4AB
`define Tile_X2Y14_Emulate_Bitstream 640'b0000000000000000110010110100010000100110001001011000000000000000001101101110000001101010010000000101010010100000000000011110000000110100100111110111100000010100001010000111000000001000010001000000000000000101010100101000000100000100000010100101100010101100111000000000100001000001101000111000000000010101110100001110010001101000000000100000000000101001101011100000000111000011100000101000110001011100010000011000011110000000000100010101001000000000000000000100011001110000001000011000000010100010011110011011000100001101111101011100100100000010000000101101011111000011000000000000000111101110110111000000000000000000000000000001010001110010
// X3Y14, RegFile
`define Tile_X3Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000001010000000010000000000000000000000110000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000011000000000000000000000000000000000000000000001000000000000000010001000100000000010000110000000000000000000000000000001010000000100000000000000000000010000000100000000000000000000000000000000000011
// X4Y14, LUT4AB
`define Tile_X4Y14_Emulate_Bitstream 640'b0000000000000000111001101000000000011111111001110011001000010000000001000011000001110100000000000110010101111000001000100000000000000000000100000110100000100010000010000000001000100000100000100001100000000111110110001100000100001110000000011100010000110000000000010001111110001100000000000000000000011010100100101101000100000000000000100000001111111000100010001000000101000000000001101000000000010000011101000000011010010000000001010000100101000101000000000001010100000000001000001001010000001001000000001011000010000000000000001101010000000000000000010111100111001000001100000000000000001000110111000010100000000000000000010011000111000000
// X5Y14, LUT4AB
`define Tile_X5Y14_Emulate_Bitstream 640'b0000000000000000010001011000100000001010000000000000010000000000000100000101010000001100010010000110010001001010100001101000000000100000000000000000000001000010011010000000001010101101010000101000000000000100010010001101001010000100000000010100000011000100111000001000010000000001100001000000000000001111100000101100101101101000000000000000000010001000000011000000000001000001000000100000100101000101000000100000101010010000000111100100000010000000000000000000000000100000000000011000000000001000000100000000000100000000000001111100000000000010000000000000101011000000001000000000000010000000000111100010000000000000100000000001000110101001
// X6Y14, LUT4AB
`define Tile_X6Y14_Emulate_Bitstream 640'b0000000000000001110000000000000000000000000000100000001010011000000001000000110001100000000110000000010100011001001001110010010001000000000111010100100100001001011010000000011010001101111100001000000000000110000000001000000000000000000000000100111001100000000000010000000010100001010001000000000000001011101000001100110000101000000001001100001111101100010001001000000010101000000000100111110100000000010101100110001010100000000011000001100010000000110000111000100010000000100000000001010001110000001000001000110011000000101001100110001010000000000000001010000000100001001000000000001011110010011110010000000000000000000000000111001000010000
// X7Y14, DSP_bot
`define Tile_X7Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000110000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000001000000000000000000000000000101000000000100000000000000000000100111000000000000000011000000000000000000000000000000
// X8Y14, LUT4AB
`define Tile_X8Y14_Emulate_Bitstream 640'b0000000000000000010000000000000000010110000000000000000000001000001001000110000000000000000000000001010000110001000000001101000000001000000000010010000000001000000000000011000010101100000000000000000010000000000000001101000100000110000010000000000011000000000000000000101000000000000001000000000000000010001001001110000000001000001101000000011100100001010010000000000010010000100000000000000000000110000100000010001000000000000010101000100100000000000000000000001010100000000000010000000000011000001001001000100100000001100101001101000000010000000000000100101101011011000000000000000010011101001011010000000000000000000000110011001000010000
// X9Y14, LUT4AB
`define Tile_X9Y14_Emulate_Bitstream 640'b0000000000000000000001100000000000010001000001011001000000011000000101000010000100100101000000100000100000000000011000000000010000001001100000100000000000010100001000000000010110101001000100100001001000000101110100011110000100001010000000000001000000000000000000000000000100011000011001110001000000010000011111001111001000100000000001011000000000110001100001001000000011010011001001001111100000001000001010000110101010000100000000100000000000010000100000000000001000010000001000001000000001001100000101000000100000000000000010001100100000000010000000010010011010000010011000000000000010000100011000001000000000000000000000000000000011100000
// X10Y14, RAM_IO
`define Tile_X10Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000
// X0Y15, W_IO
`define Tile_X0Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001100100000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y15, LUT4AB
`define Tile_X1Y15_Emulate_Bitstream 640'b0000000100000000001010000000000000000001100001110000000010001000000100000011000111101001000000000000010010010101001101000010000000100000100000110010100001100010000000000010001011101000100000100001011100000110010100001110001100001100000000100100001011111000000000000001101100100000100010000000000000010111000100101111110000001000000000000001000011000000000010000000000101101000000000001100010000100111001010010000010100000000000011000000010000000000000000000001001000000000001000000000010000000101001010010010110000000000000010001000000010000000000000000001100100100000000100000000000000110001010100010000000000000000100000000001100100000000
// X2Y15, LUT4AB
`define Tile_X2Y15_Emulate_Bitstream 640'b0000000000000000010000010000000000000000000000000000000011000000000100000001000000000000000000100000010000000001001101000100000001100001100000000101000100000110010010100100001001000001001000100001000100000001000010011010000101011110000000100001010011001010000000010001101011000000101001010011000000010000101110000000001000000000001010000000000110011101000000001000000110110100100001000110000100010001111100001010000000001100000001000101110000010000000000000010000111000100000111010000011000001000000011100011000100000000000000000100100000010010000100010001011000000010001000000100001000000000000110110010000000000000000000000001000101011010
// X3Y15, RegFile
`define Tile_X3Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000000100000000000000000000111100100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000010000000000000000000000000000000000000000000000000000001000000010000000110110011100000000001101000000000000000000000000000000000000000000000000000010000000000000000011000000000000000000010000000011
// X4Y15, LUT4AB
`define Tile_X4Y15_Emulate_Bitstream 640'b0000000000100000000000001001000000000110000000110110000000000000000001001011000101111100000110000111000111001001001001100110010000000101000111000001100100000011000010000100110010101100011000000000000100000101000000000101100000000000000000110000110001000000110000000000010000101100001010111000000000001110000010000000000110101000000000010010000011111000011010000001100000000110100001100000110000000000000010000000001010000000110010110000000100100001000000000000000000110000000000001000000001110000000100000011000100000000000110010000000000010010000000011000011011100000001000000000101000100001100001001000000000000000000000001000000010000010
// X5Y15, LUT4AB
`define Tile_X5Y15_Emulate_Bitstream 640'b0000000000000100100001001100100000001000000000000000000000000000000000001100100111101000101100000000000110000111001001100000010001000100000100000001100000000011011110000000000100000000000010000001100000000000000001000001001000001000000010001000000001000000110000000001110001000000000000000000000000000010001010011100000000111000000010001000011000011100000101000000000000011001000001000000110000010000110100000000000101000000000000000000000010000000000000000001000001000000000000000000100000001110100000000000000000000010000100000111100000000000000000011011100100010010000000000000000110010010010110001000000000000000000000000000000000011000
// X6Y15, LUT4AB
`define Tile_X6Y15_Emulate_Bitstream 640'b0000000000000100100001001110000000010100111000000000000000101000000101100111000100001100000010000110000001100100000000000000000000100001100011110001110100000000011000000010110010100001100110101001000000000010000100011101010100001000000000101101000011010000110000000000010010100010000000010000000000001000100001001111000110111000001001111100000011000001010011001000000010000010000000100110100000000001010000101000000000000100000000011000000000000001000000000100001000100000100000000000000000000100011000001000000100000100000011000010010000010000000000110001001000000011010000000000000000000001010001011000000000000000100000000001000010010000
// X7Y15, DSP_top
`define Tile_X7Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000001100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y15, LUT4AB
`define Tile_X8Y15_Emulate_Bitstream 640'b0000000000000010100000110000000000000000101000001111000000000000001100100000000100010000110110000000100000000110010000100010000000000000000000011010100000000000001010000001101100101101000010101001100000000000100011101101001111011000000000000000101011001011000000000000001000000000100011000000000000000000000010000011001101101100000000101000000011000000000001100000000000000011000000000110100001010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000010100011000000100000010010000000010010000010000011001100000000000100000101101000000010100000000000000000000000001110101000
// X9Y15, LUT4AB
`define Tile_X9Y15_Emulate_Bitstream 640'b0000000000000000101010111101000000100000000000111001010001000000000000000000000010110000010100000001010000100000000000000100000000011000100000000111100000000000010100000000000000100000110010000001000110000000000000001100010000001100000010000000100001101000000000000000000100000000011010000010000000000001000101011100000110001000000100000100010000110101010110000000000001100010000001000111000000000010000000000000001101000000000001010000000000000001100000000001110000100000000000010000000000100010000000001011000100000000000011000000000000010010000000001101001000000000000000000000001100011101000110110010010000000000000000001000111101000000
// X10Y15, RAM_IO
`define Tile_X10Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000
// X0Y16, W_IO
`define Tile_X0Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y16, LUT4AB
`define Tile_X1Y16_Emulate_Bitstream 640'b0000000000000000000000001100000000000000000000000000111011001000000100000000000100000000110100000100000000000100000001000000010001000000000101101101000000000000000010000000001110000000000010000000110010000000000000100000001000000000000000011000000001100000000000000000000000110000000000000010000000000001010010000100010100000000000100000001000000110000000000000000000001001110100001000000001010000000000100000000011000000000000010000000000000100000000000000000000000100000000000000000110001000000011100000001010000000010000000000000100000010000000000010101000000000000000100000100000101000100010000001000000000000000100000000000000000010000
// X2Y16, LUT4AB
`define Tile_X2Y16_Emulate_Bitstream 640'b0000000000000010100100001000000000001011010001010000000000000000000001100000000000000101110110000110000100010000010001110010000000100001100000111111110001000000000110000000011010101000010110100000100000000001110100100100010000000010000000001100001000101000110000001000001000100000011000000000000000100010010000001000011000010000000000100000000111000001000000100000000100000010000010000110001000000110000011011000010110000000000011010001000000011000000000011000010011110000000100011000000000000000001000001011010100000010010100100000100000000000000100010011010101000110010000001000001000110001010000011000000000000001100000010000101010010000
// X3Y16, RegFile
`define Tile_X3Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100100000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001010000000001010010000001100000000000000110000000000000011000000000000000000000000000000000000000000000011000000000000000000000000000000000
// X4Y16, LUT4AB
`define Tile_X4Y16_Emulate_Bitstream 640'b0000000000000001000001010000000000011100000001110011110011001000000000100001010001110011011110000000000000001001001000000000010001010000000000010000010001000000000110000100000000000000000000000001000100000101000110000000000000001110000000100001000000101101000000000000100000000000000110000000000000001100000100000010000000001011000000000000000010100000010000000000000100000000000000000111001000100000000000010001000000011000000000001100000000000000100000100000000110000000001100000000010001100000010000001010010100000000000000100000001100010010000000010010000000000000001100000000001100000000110000000000100000000000000000001000000000000000
// X5Y16, LUT4AB
`define Tile_X5Y16_Emulate_Bitstream 640'b0000000000000101100001001100000000010100000000000110000000000000000000000010000000000101000000000001000000101000110000100010000000000000000011001000100100001011010000000100100001100001010110100001001000000101000100000101010101011000000000110000010010001000000000000000011000111001001011000000000000000110000100000011100100101001000001001010011000100001010011000000000000000001000000000110110001000100010000001000011000000000000111101000100100000001000000000000001000100000001100000001000000000100011000000000000010000000000000000011100110000010000000000000000010000010000000000000000100011000000000001010010000000000000000000000000000000001
// X6Y16, LUT4AB
`define Tile_X6Y16_Emulate_Bitstream 640'b0000000000000000011000010000000000000000011000000000000001111000000001100000000000000000000000100000000000000000010000000000000000000000000000000000000000010010000011000010000001000000010000000000000001100010000000101000000000000000001000000000000001000100000000001000000010000000000000000010000000000000000000100000010000000100001000001000000000010100000100000000000000000111000001000001000000000000010000010001000101000000000001010100000000000000100000000000010000000000010000000000100000010000000100000000000000000000000000100001000000000000000000011100000000011011000000000000001110000000000000010000000000000000000000000000000111010000
// X7Y16, DSP_bot
`define Tile_X7Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000
// X8Y16, LUT4AB
`define Tile_X8Y16_Emulate_Bitstream 640'b0000000000000000011000010000000000000000000001000000000000000000000000110101010100000000000000000001000000000111001000000000000000010000100000011010000000000000001000000100001100100000000010100001000100000001000000111100000100001000000010001100000101000000000000000000000000000110000011010000000100000000010101001100110000100000000000111000000111101100000001000000000000100010000000100000100000011011001000010000001000000000000010000001000010000000000000000001100000000000001000000000000000110000000000100010000000000010001101001100000110010000000000000000000011100000000000000000000010011000000000010000000000000000000000001010000001000000
// X9Y16, LUT4AB
`define Tile_X9Y16_Emulate_Bitstream 640'b0000000000000001101000100000010000100000000000000000000000000000000100000011100011000001100000000000110010010001001000000000000000001001100000110110000000110010000000000010000001100000111111100001110010001010010000001000010100001110000010000100000101101000000000000000100001100001010011011011000000000001001111000000001010001000000110000000011100100000111000000000000001011000000000001110000000010001100000000000011110000000000001110000100010000001000000000000010000100000000000001000000001001000000000001000000000000001000111000111000000010010000000000100011010110000000100000000000100101101000000010000000000000000000000000001000011100000
// X10Y16, RAM_IO
`define Tile_X10Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
