library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package emulate_bitstream is
--X0Y1, W_IO
constant Tile_X0Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y1, LUT4AB
constant Tile_X1Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X2Y1, LUT4AB
constant Tile_X2Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X3Y1, RegFile
constant Tile_X3Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y1, LUT4AB
constant Tile_X4Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X5Y1, LUT4AB
constant Tile_X5Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X6Y1, LUT4AB
constant Tile_X6Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y1, DSP_top
constant Tile_X7Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X8Y1, LUT4AB
constant Tile_X8Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X9Y1, LUT4AB
constant Tile_X9Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X10Y1, RAM_IO
constant Tile_X10Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y2, W_IO
constant Tile_X0Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y2, LUT4AB
constant Tile_X1Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X2Y2, LUT4AB
constant Tile_X2Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X3Y2, RegFile
constant Tile_X3Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y2, LUT4AB
constant Tile_X4Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X5Y2, LUT4AB
constant Tile_X5Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X6Y2, LUT4AB
constant Tile_X6Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000";
--X7Y2, DSP_bot
constant Tile_X7Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X8Y2, LUT4AB
constant Tile_X8Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001001000000000000000000000000000010000000000000000000000000000001100000000000000000000000000000010000000000000000000000000000000000000000000000000100000100000000000100000000000000000000000000010000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X9Y2, LUT4AB
constant Tile_X9Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X10Y2, RAM_IO
constant Tile_X10Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y3, W_IO
constant Tile_X0Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y3, LUT4AB
constant Tile_X1Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000100000000000111001000000000000000000000000100111110000000000000000000000001110000000000000000000000000000000001100000000000000000000000000001000100000000000000000000000000000100000000100000100000001000000001000000000000001000000010000000001000001000100000000000010001100010000000000000100000100000000100000000000000000000000000000000000001010100000000000000100000000000000000000000000000001000000001000000000000000000000000000000000100000000100000100000000000100000000000000000000000000100011000000000000000000000000000000000111000000000000000000000000000000000010000000000000000000000000000000000000000000";
--X2Y3, LUT4AB
constant Tile_X2Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100001000000000000100000001000110000000000110000000000000000000010000010000010100000000000000000000000000011010000011000000000000110110010110011001100000001000000001101100000100001110100000000000000000010101100001010000010000000000000001001001000000000000100000000001010000010000000000000001100000000100101101000000100001010001100000101100001010000000000110000000000001111111000010101000000010110000000000000000011000000100000010001100000000001000000100011010000000000000000001001100100101000000000000000100000100110111000000000000000010010000000101000100000000000000100000100000001000010000000000000000000000000000000010000";
--X3Y3, RegFile
constant Tile_X3Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y3, LUT4AB
constant Tile_X4Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000011101000000000000111110000000000000010010101000000000010000000000000000010010000000000000000000000100000111000000100000000000000100010011000000000000000000001010101100011000000000000010000000000110000100100100000100000000000100001010101000000000000000000000000001000000001000000000001101000000000011000010000000000100001000001100000000001000000000000000000001000000000000000100000100000010000000000000100000000011010100000000000001000000000000010000100000000000000000000001000101010100000000010100000000000010100110000000000000000000001100011100101000000100000000000000000110101001000000000000000000000000000001011000000000";
--X5Y3, LUT4AB
constant Tile_X5Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000000000000100000001000000000000010100000000000100000000000000011000010000000010000000000110100011111000000001000000000000010000011000000000000000000000100000000110000100001000000000000110001100000000100001110000010001100100000000001000000000000010001000110100110000000000000001110001100010000001100000100000000001010010000101000000100001000000000010011000000100110000100000111001000000000011111000100000011110000000000000000000000000000011001000000000000011000000000001001000000000000000100000011000010100000000000000000000000011011001110000000000000000000001000001000110001100000100000000000000000000000001000000000";
--X6Y3, LUT4AB
constant Tile_X6Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000001110000000000000001010101000000000000000000000001000110101000110000000000000100001100001000110100000000000000000000000000000011010000000010011000001000101101000000001000101101001000000001010010000000001001110001000000000100100000010010001001000010000000000100111000000011000000000001101000100000000000001100000000001101000001100000000001000000000000001100111000000000111100000010110010000000000000000000000000011000001000000000000110000000000010000000000000000000000000000000000011100000000000001000010000000100011100000000000000000001011011000001000000000000000000010000001000000100010000000000000100000010001100000010000";
--X7Y3, DSP_top
constant Tile_X7Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001100000011000000000000000000000010110000000000000000000000000000000000001011000000000000000000000000000000000000";
--X8Y3, LUT4AB
constant Tile_X8Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000010100001000000000000100111100000100000000001110000001000010000100011110000000110000011100000001010100000000000010000001001000000000010000000001001000000000101000000100000001100001000000000000100110000000100000011010110000000101101000100101010000000000001100011000000010011110000000000010000101010000000000100000000001000011110000011110000000000000000000000110110100001000110000000000000001000000000001000000000000000000100000110000000000000000000000000000000100000010000000001001011100000000000110000000000000110000000100001000010000000010101001010000011001000000000000101010000101000000000000000000000000000000000000000000000";
--X9Y3, LUT4AB
constant Tile_X9Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100001000000000000000000000000000000001010011000000000000000000110000000001000000001100000000100010000000000010000001001100011101100000011000000000000000010111110100000000010100001000000001010000000000000010101011010000010000000000000000110001000000001100010000000000001000000000000000000011100000000000011000000001001000000000000000000010000000000000000010000000000000000000000010001000000001000000000000000000001000000000000000000000000000000000000000000000000000000000001001000001100000000000000000000000000000000000000010010000000000100011000000010000100000000001100000000100000000000000000000000000000000000000000000000";
--X10Y3, RAM_IO
constant Tile_X10Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000";
--X0Y4, W_IO
constant Tile_X0Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y4, LUT4AB
constant Tile_X1Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000100100000000000000000010001000000000110010010101000000000000100000000000000000000000100010000000001001001000000000000100101100000110100000010000011000000000010011010101100001100000000000000001010110000001100100001010100000010000000000000011010110010000000100101000010101011001011100000000000000000000011000000100000000000011000000100011001001000001000000001001000100001000110100000010000000110000000000100001000000001001000000011000000000000000000000000000000001000000000000000000100000001010011100000000000100100000100100010000000000010001011101100000111001000000000001100000001001010100010000000000000000000000000000001000000";
--X2Y4, LUT4AB
constant Tile_X2Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100001000001000000100000001000000000111001110000000100000000000000001111111000000001110000000000110100001001010000001000000001100010010000000000000000000100000100001100000011000000000010001001000100001001010000000110000000000000000001000100001000000001100001100000000000111010000000000000001000001000000011000000000100100000000000110000011000000000000000011000000001000000000000000000000100000000011100001000000001100000001010000000000000000000000000100000000000000000000000000000001101001011100000000010000000000100000000000010000000001001011000100000001000000000001100011111000000010000000000000000000000000000000011000000";
--X3Y4, RegFile
constant Tile_X3Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y4, LUT4AB
constant Tile_X4Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000100000101010000000100000001001010000001000011101010110011100011110100001000110000001000000001000010000101000000011100010010001010010000000000100110011100101000110001000000000100001110100001101010010000101000000001100000001010001000000001001110101100000100000000010000010011110000000101100110110010000000110000000011100111100010110000010000100000000010001000001010000000000101000110001111101000000000000100000000000000000100100000001000001000000000000000000000001000000100000000000100000000011000100100011100000010000000000000000101111000000000000000000000001110000101111010010100000000000000000000001000100011001";
--X5Y4, LUT4AB
constant Tile_X5Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000110110000000000000000000000000000000001010110000000000000000000110001010000000000000000000000000110100001001000000001000000000001010010010000010000000000011000101001100000000000000000000000011110000000100000001010110000000010001000000000010000000000001001110000000110001000000000000000100111100000000001000000000001001001000010011111001000000101000000101010011000001100110000000010101000000000000001010000100000000000010000000000000000000000000000100000000000000011000000001001000000000000000000000000010100110000110100000000010000000010110000100111010000000000001001001010000000110000000100000000000100000100001100000000000";
--X6Y4, LUT4AB
constant Tile_X6Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000010001100000000001000000011111010001111000000000001000000000000000010011101100000000000010000111000011101001101010000001000001000011100011100000000010010010100001111001101100011010000000100000000000000001110101111000000000000010000000100010110001001000000000001101000000001000111001000000000001001100100011000101010000000010011000001100000101001000000000000000000000100000000000010000010001100010000000110000100000000011101000000000000000110000100000000000000000000000000000010000000100011100100011000000000001000100000000101100010000000000011100110000000011010100000001000000000000000000100001000000000000000000111000011011010000";
--X7Y4, DSP_bot
constant Tile_X7Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000111000000000000000000000000000000100000010000100000000000000000000000000111000000000000000000000000000001110010000000000000000011000000000000000000000000000000";
--X8Y4, LUT4AB
constant Tile_X8Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000110101000001000000100101010001100110011010111000000001100111010001010001001000000001100000010001011100000010010000010001000000110100100010001010000010000100101000001100110111101000110100000000000101001001000010000000000010000000010000100000000000010000001100001000000000011000000000000000000000101011000110010000000100101000000011101000011010000000000001000101000001100001000000000100000010011000111010000100000000000001000100000001100000000000000000100000000000001000000001000000010100001000010001000000100110000100100000000000000000011001000010000010000100000000000111011101001011000000000000000000111000000111000000010000";
--X9Y4, LUT4AB
constant Tile_X9Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001000000010000000110011000001011111011010000001101110011100010000010110100000011100001000000000000000110010000001001100000000011110000010011000010000000100100001100000001100001100000100000000000001000000100001010000000000000010001100010000000001000000001000000001000011000000000000000001100000000000000110000000011010000000000000001001001000000000000010001000000000000110000000000110100000000000000000000000000000000000000000000000000000000000000000000000000010000000001101000000100000000010100000010000001010100100000000000000000001000000000000000000000000000000000000001000001010010100000000000000000000000000000010000";
--X10Y4, RAM_IO
constant Tile_X10Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y5, W_IO
constant Tile_X0Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000011000001100000000000000000000000";
--X1Y5, LUT4AB
constant Tile_X1Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000111000000000001100000000000001010101001011001000010001000001000111000100000100011000000100010000100000010010000000110000000110000000000000000000001000100000000000010001110001101001110000000001100101000010010001000100000000100000010000100000001000100000000001000100101000100000111101000001100000000000001000000001100000000001100100000000011110000101000000000000000001010010101001001000000010000001001010010001000000000000000000000000000000000100000000001001100000000000010010000000001000000001100001000000100000000000001100000100000010000000000001001001000000001000100000000101100010001010000110010000000000000000100000000001000101000";
--X2Y5, LUT4AB
constant Tile_X2Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000010000000010000000000011110000001111111000001010000001000011000010010011100000110100001100000000010100000101000010001100100000001000011110000010111010010000100001010000000000100000000110000100001110110000000001000000000000000110101100000100000110000000001111111000000011110100011001100011110001010001111001100100000001110011000001000110000100100001000000100011000100001001001100000000000100000000000101111000010000001111000000000000000100000000000010000110000000000001000000001010000000001001000100100000000100010101100000010000000000000000000000000000000000000000000001111010111011010000000000000000000000000000001001001000000";
--X3Y5, RegFile
constant Tile_X3Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000111000000000000000000000000000000000000000000000000";
--X4Y5, LUT4AB
constant Tile_X4Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000010000001100000000011111111000101100111001110000001000011000010010011100010110100001000100000010100000001001010000000101000111000100000000011100000010000101111000001100001111001000000010000111010001100000101011010010000000100101000000000011111000000001000000101000000001111010000000011101000001000011000001000000000000001001100100110100001010000000000101000000000001000001010000010100000000001000001000000000000011111000000000000000000000000000010000000000000101000000000001000000011100101000000000000000000000000100101000000000000000001111111001100011000000000000001101010010010010111000000000000000000000101000001100010000";
--X5Y5, LUT4AB
constant Tile_X5Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000011100111100100000001010101000000011010010101000001000111101000010010011010010000001000110001110100000011001000000000000000011111110010011000000000100000101111110101101000001001001000010000111110100001101000010001100000000110000100001000000000000000100001100101000000001000000000000000100010101110000001000011000000110011000010000111000000011000000000001100010000001100000010000010100101000000000001010000000100000100000000000000000000000000000000000100001000000001000000001000000000000000001000000000000100111000000100000000010000000001111100101000000001000000000000101101100010000011010000000000000110000100001101010010000";
--X6Y5, LUT4AB
constant Tile_X6Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000100000000110001000000000000101000100001100000001001110000000000010100010011000100111110000001110000000011101000000011010000011101100011110110000000000000011010000011111000000000000010000000100100001010010101101000001001010010000010000000100001101010110000000001100010000000101111000011000000000001001110010000000100100000001010101000011100001001000101000000000010100100000000000111100000010110101000010000000001011000000011010100100100000000100000100000001000100000001100000000010001000010111000000011010000000001100000100111100010000000000000001001010000101011000000000000000101000000100110100010000000000000100000110110001111001001";
--X7Y5, DSP_top
constant Tile_X7Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001100000000000000000000100000000000000000000000000000000000000000000000000000000010100000000000000000000010100000000000000000111100001111000000000000000000000000000010100000000000000000000000000000000000000000000000000000";
--X8Y5, LUT4AB
constant Tile_X8Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000100100100000001000000011111010000000100101000101000001101000011000110000000101010000110000111010010110100000000000001110000000101000011000000000100010100100000000110100001100110000001110100000100010000000101111010001100000000010100000010100000110000000000010101100000100000100011000000001100011010001111000110011000000110000000000000100000110011000000000000010000100001001001000000000010100111010000011100000000000000010010000000000000100000000001000010100001000000000000000000001110010001000000110000000010100000110100000000010010000000000010001111001000001000000000000100101101010111110000000000000000000000000001100100010000";
--X9Y5, LUT4AB
constant Tile_X9Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000010000000001000000001001100001111000111010000000000000001000010001100101000000000000000011010001001000010111000000000101000111100000000010001000000010000111110000001100001110001000100000000111110100001010100010000000000000110000100000010100111000100000001100000000000000101000000000000100000000011100000001000000100000000010010000001000001000000000011001000000100000100110000000000100000000000100000110000000000000110000100000000000000000000000100000000000000000001000000000100000000100001000000100000001001110010000100000010010000000011100001100100000001100000000000110000000000000100010100000000000100000000001001000000000";
--X10Y5, RAM_IO
constant Tile_X10Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000";
--X0Y6, W_IO
constant Tile_X0Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000010100000000000000000000000000011100001110111000000000000000000";
--X1Y6, LUT4AB
constant Tile_X1Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000100001111110000000000000000110011000010001000000001000001100110000100000100011000000100101100000000000000100000011000000111000100000100000010000010000000000000000001000001100001010000000000100000010000101010000000000000110000000001100000000001000100000010000000001010000100110000011001100000010011100001111010100000000000001000000000000000100000100000000000000010000100000100111010000000000100010010000000001000000000011000001000000000000100000000000100000100000100100000000000000100100100000000000100000000001000000001100001000000010000000000001100000100000001000000000110010000000101000000000100000000000000101000000100000100000";
--X2Y6, LUT4AB
constant Tile_X2Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000010000000000000000000000011111111001100010000001100000001101110011010001000101001110000011110001001001101100100011010000011101100000001100100111000010000110000010101111100000000001000000000100000010110100000100000000000010000000101100110000001000110000000000000111001000001010011011000000000000011011001111000000000000000010000000001101100101001110000000100000010000000000000111000000000000101000010000001100000000100000110100100000000000100000000001010001100000000000000000000001000000100001000000000000000000000100000011100000000010000000001000000100000000000000000000001110001001110001000000000000000000000000000001000010010000";
--X3Y6, RegFile
constant Tile_X3Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000";
--X4Y6, LUT4AB
constant Tile_X4Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000010000000000000000000000011000011001011111001000010000001001100100000100110011001000000000000000100000001000011111010000001000000000000000100000001100000000000100000001000000000110101000101000000010110100011100010011010000000000110101000110000000000000000000010001000000001101110000000000011100100101010010000010000000000000000000011100110000110011000000000110100000100001001000000000010000001000000000001000000000000000000000000100001000000000000001000000010000000000010000000000000000000000100000100100000000000110000110100000010000000000001010111010000010001000000000001101101000011001000010000000000000000000000000001000010001";
--X5Y6, LUT4AB
constant Tile_X5Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000011000000011000110001111000000000000000000001000100000011110000010000000000000100101010001000000000000000000000000000010100000000000010000000000100000001101101010000000000000000001001110000011100000100000100000010001100000100111001000000000001111011000011100111110011000000001100010101010011000010000000001011011000011100000100010100001000000000001000110000000110000000010000100110000010000101000000110000010000000000000001000000000000001001000000000000000000000001000101100001100001100000000001000010000011000000000000000000011000011010001000000100000000000001110010100000000000100000000000000000000000001000000000";
--X6Y6, LUT4AB
constant Tile_X6Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000100111101100001000000000110101000100111100011100000000000111011110011010100100110000000010000001100010001010110000001011000000001011111100001101000000000100110000101100000100100001000010110001010110000000100000011010010000010011100110010000110001000000000101011000000000001100000000000011100001000011111000001000100001000001001110010011100100111000000000000010000000000001001000000000110010000101000000101000000000010000000000000000000100000000000000001010000000001010000000001001101101101000011100100000000000100010100100000000010000000011000011110100010001000000010000111110010010001000000000000000000000000000000110001000000";
--X7Y6, DSP_bot
constant Tile_X7Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000100000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X8Y6, LUT4AB
constant Tile_X8Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001101100000000000000000000111111000010010000000000000000000111110100000000100100000010000010100000111110010001100000000011101111100010010010000000000000001010100000000110100001100001000000000001001100000100001000001010000000100001000000110000000000000001000000100000000011000000000000010100001000000000000000000010100000000011010000000000001000000000000000000001000001010000010000100000000000100000000100000000100000000010000000100000000000000000000000001001000000000000000000001101010000010000000010000101000000000010010000000000000010001001000000000100000000001101010000111001000000100000000000000000001000000001100000";
--X9Y6, LUT4AB
constant Tile_X9Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000100100000000000100000000001111111101010000000000001110011010000010010101110000001010000000000010100000110010001000100000011101101110001100000010010000001111010000000101101000000100010000000000000000000000000000110000000010000000100001000110000000000001001000000000010011010000000000100011000000000000000010000000110000000000000011000101000000000000000010000000001101010010000000100100000000000000010001000000001010000000010000100000000000000000000100000000001001000000000011000000011001000000000000001100110010100000000010000000000001100000100100100000100000000001101001101100110000000000000000000000000000110111000000000";
--X10Y6, RAM_IO
constant Tile_X10Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000";
--X0Y7, W_IO
constant Tile_X0Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000001000000000100000000000000000000000000000001011100001110000000000000000000000";
--X1Y7, LUT4AB
constant Tile_X1Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000001000000000000100101100010000000010011000010000001010110000000000111001000000000000000000000000100000000000000000100100000001011100100001100110100000111100001000000111001000000000101100001000110100001000110000000000100110000110000010100000100010101000000000010000100100100000110000101000000100100000001101000000001100100000000101011010011100101100101111001000000001111000000001100001110110000100011100010000001111010100001001001001000101000000100000000000001000100000011100011000100001001000000001011011010101000001100000000000100010010000000000001101111010000001000100000000000001101110011100000000000000000000111001001110001101000010";
--X2Y7, LUT4AB
constant Tile_X2Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000010000000000010000000000000000000000010001010000000000001000111000000001101001000000110000001000000000000001011000000111001000000000001010001001000000000000000010001001100001110001000000100000111000000101000100010000000000000000000010001000000110000100001000010000000010000101000010000100000100000101000100000000000000000101000100000000001000001001000000110000011000000000001010000010000010000011000000000000001000000110100100100000000101000000000000001110000101000010010000000011001000000001010010100000000000000100100100100000000000000000100000000100000001000000000000000000000000001010000000000000000000000000000000100010001";
--X3Y7, RegFile
constant Tile_X3Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110000000000000000000000000000000000000000000000000000";
--X4Y7, LUT4AB
constant Tile_X4Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000010110001000100000000101001110000100111000000000000000101000110010000010011000100000010110110110000110100000111000000000000000000010011110000001000001100000010000100000001010110001001000000000111000101101010001010001010000000100100000001010100001000010001000011000010010010000010000000001001000110001111011111101000001000011000000000010101000011000000000100101000000001000010100000010001000000100000000010000000000001010000000000000001000000000001000000000000000001010000000001000000000100100000000101000010100001000010101000000010000000000000001001011001000000000000001110000000011001001000000000000000000000000110000100000000";
--X5Y7, LUT4AB
constant Tile_X5Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000001101001001000000000000010011001001011011110011101000000100100001100000100000000000000010100110110000001000000110000000001101100000100001000011001000010010000100010010000000000100001000000010001001000000001000000010000100000010000000110000100000110000000001100001000001001000000000000000010000000000000000110000010000000110100000010000000100000100100000000110001000000000000000010000010001100000100000000101000000000000010000011000000000001100000000000000100000000100000011000001001000000101001011010010000001000101000000100000000000000000000100010111000001000000000000000000000100000000000000010000000000000000000000000010000000";
--X6Y7, LUT4AB
constant Tile_X6Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000100000010000001000000000000001100000000011001000010000001100010000000010010011001000000100000110010000100000000110010000100000000000010010000001001010000000000001000111101100110011000000001011000110010000101100000101010101001000000101010001000110110000000001101110000011000011000000001110010011100000000000000010000000001100001010000000110000010000000000000001000010000100000000000000010001011001001010000100000000000000000000000000000001000000000011001010110001001100000000001000010100000000001000000000000000000000011100100000010000000000000000001000000010000000000000000011000100000001110000000000000000000100001000000000100000";
--X7Y7, DSP_top
constant Tile_X7Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001100000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000011010000000000000000000000000000110100000000000000000000000000000000";
--X8Y7, LUT4AB
constant Tile_X8Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000101010000110000000000100001010001000001111011010000000000110000010000010000011000000000010001000001101001000000010000001000000000010110000101000000000010000100001101001101000000101001110110000001100000001011110111011000000010010101010001011011000000000000011111000000000011000011000000000010100100001100000100000000001110000001000000011000000001000000000000000000110001000110000000010001100000101000010100000000000001001000011010000000000000000001000000110010000100010000000000001100010100000000100100000011000001011111100110000000000000010000011000000110000100000000000100000100000001000010000000000000000000000001000000011010";
--X9Y7, LUT4AB
constant Tile_X9Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001000000000000111110101000000011000000000000000000110000000000011111010000000001110000001000110100001111010000010101100011110010000001000000000010000100110110001100001010100001001100000011000000000000110100011101000000000001000000000000110000000001000010010001100000001010000010010000100100010011110010001000000000000010000000100000011010000010000100000000000000000001000000011011000000000000011100000000000001101101000000000000100100000000011000000000000000000000000000010100001100000010000000000010000000000100000000000010000000011000011000100000000000000000000001011010000000000000000000000000000000000000001000000000";
--X10Y7, RAM_IO
constant Tile_X10Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000011000000000000000000000000000000001100000000000000001000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000010000000";
--X0Y8, W_IO
constant Tile_X0Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001110001000000000100000100000000000000000000000000111100001110000000000000000000000";
--X1Y8, LUT4AB
constant Tile_X1Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000001000010000010010110000110000000000000001111001000000100000001101000000000000010011000000000011000001000010110000000011000001111101000000001000000000110100011000100000100000000001111000000000110100000000000010100000101001010100000010001000100010101010000000000001100000010000100011000010000000001000001010001100010000001000000100111000000111001000000001000000000000011000100000001111100000010000001100010010000000000000000010101111001001000000110000000001000010111000000000010000000010000000101110001001110100001000100000000100000000010000000000000010011000000010000100001010111100000100001100000000010000000000000001001011100010000000";
--X2Y8, LUT4AB
constant Tile_X2Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000110010000010000000001000100001010000000000001000000000010001000000100010000000000010100010000010001101101010000000001100000000100001100000000000000000010101001000101000000001000000010000000001010000001100001000000100110010000100100001100001001000000000000001000000000000111011001101001101000000101100000011000000000010100001110011100000001011000000000001000010100000000000000100010100100000011000000000011000000010000010000101000000000000000000001000010000001000000000000001001101111100010010000001000010100001000000000100000000100000001100010000000000000000000000010101101001000100110010100000000000000001001001010000001000";
--X3Y8, RegFile
constant Tile_X3Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y8, LUT4AB
constant Tile_X4Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000010000000000000100000101010101001111000000000111000001001000010000001100000000000000010000110110000000100000000010000011100000000000000000010001110000010000000001011100000001111001000000100000011000001010101000011010110000000000000000000000110110000001000000010101000000001100010000100000000011000100011111000000000000000000000000010010100100111000000000110010000000001001011000000000000010110010001000101000000000001010001001110000000100000000001000000000010000000000000000000001111100000010000000000000001000100000100100100000000000000000010011110000110000000000000001101010011010001000010100000000000000010000110011000001000";
--X5Y8, LUT4AB
constant Tile_X5Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000011000000000000000001010101001001001000000011000000000000000100000000000000000100000010000000000001100000000000000000000000100000010000000011100001000000001000000101100000110101001000000101001010000000110010110001000000000000100000000010000000010000000100001001000000100100011000000010000000101000011000110100000000011101000001101100000110111000000000000000101100000001111100000010101101000111000001001000000000010000000000110000000100000100010000000010000001000000000000001001100000000000000000000000011000010001100100100000000000000010000101010101001000000000000001100011000100010100010000000000000000000100001000000000000";
--X6Y8, LUT4AB
constant Tile_X6Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000001111000000000000000101001100001110000000000001000001001101111010000000000000000000100000000010000100000011110000001100000000000010110000000000011011100000001001010001101010000101001000010000110010000001001000110001100000000000001100000100000110000000001100010000100010110100000000000010001101100001100000110101000001100001100000111001000010101000000000000000011000000100000110000010110000000111000000011000000000010110100000100000001000000000000010000000000100000001000000011000000000000011000000100001001000000101100100010000010000000010000101010100001000000000000001010000100100111000000000000000000100000000000000000000000";
--X7Y8, DSP_bot
constant Tile_X7Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000110001101000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000100000000000000000001000100000000000000000000000000000000000000000000000000000000000000100000000000000000011000000000000000000000000000000";
--X8Y8, LUT4AB
constant Tile_X8Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000010000000110100000000111110000000001111000001111000001101101011000000010000000110000000010011110010110100000000010000000001000100000100000010000100000000000110010110000000111100100001000000001000110000000000100100001000000010110000000000000010000000001000001100000000010000101000000000000100000100100011101010000000000100100000000011110000011001000000000000000010101001001000000100000001000010010000001010000000000000000000000000000001000000000000000000000000001000011100000001000100000000011001000100000011000000100000100000000000000000000100001011001001001100000000001100111100000000000000000000000000000000000000000100010000";
--X9Y8, LUT4AB
constant Tile_X9Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000100000001010000100000000000000001111111010010101000000100000000010000010000010010000000100010000000000100000000000000000001100010100000000011000100000000000010110110100000000010100001000000000100000000000010010100001000000000100000000000110000000000001000000000000001001000100000000000000000010100000011100010000000001000000010001100010001110000000000100000000010000001001110000010000000000010000000000100000000100000000000000000000000000000000000001000000000000000000000000001000100011000000011010000000010000000011010100000010000000000000100111000101000000100001100001100101000000000000000000000000000000000000100000000000000";
--X10Y8, RAM_IO
constant Tile_X10Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000110101000000000100000000000000000001110000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011";
--X0Y9, W_IO
constant Tile_X0Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000111100001000000000000000000010000000000000000000000000000011100001110000000000000000000000";
--X1Y9, LUT4AB
constant Tile_X1Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000100000010100000000000000000000000011001111011010010111000001000001000000000000001000000000000000001000010110000000010000000010000000100000000000010000011000010000001001000101000110100000000100110000000010000000110011001010100000000000100101000011110001000000000000101010001000101000011000000000001100010001111000111101000000110001000010000000000010100000000000001000000000000100111100000000000111000000000010101000000000000111011010000010001100000000000100011100000100000000000000001010101100010001000010000000000010000001100000000010010000000010000001101111010000100000000100110000111001001000000100000000000001000001010001100000000";
--X2Y9, LUT4AB
constant Tile_X2Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000110101000000001100100000000010011000000000000000010000000000010001001000000000000000001000000000000000000001011100000100000010000001101000010010000000000000100000110101001000100110101010000000000100000010000100000000100000010000000000110000000000000000001000100000111000000000000000001000000011100010000000000100000000011111110100111110000000000001000010000001101001000000011110000010010000000101000000000000111101000100000001100000000000110000000000000000000001000000000100110100010011010100000001010100010111000100000010000000011011101100101001001100000000000000101110110111001000010000000000000000001000011001110000";
--X3Y9, RegFile
constant Tile_X3Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000111000000000000000011000000000000000000000000000000";
--X4Y9, LUT4AB
constant Tile_X4Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000011000100000100000000001110000001111011101001111000000000000010000001010100000010000000000000001000000000000000000000000100000000000000000010000000000010000100000010100101010000000000010000000000000101101110000000000100000000100100000000010000110000100000000000111000110000000010000000011001000011001101011000000000000000000001101000010100000010001000000100000000000000000010000000000000000100000110100010000100000010010000000010000000001010000010000000000000001000001000000001000000000001100000000000000000000010000000000000000010000000000100010010000000000000000000000010000011000001101000100000000000000000000110101000000000";
--X5Y9, LUT4AB
constant Tile_X5Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000010010100011111000100000000000000000001010000010010101000000000000000000100100000000000000001100000000100001000000000000000000101000001100000000000000100000010000000000100000000000010000000000000001000000001110000000001010000000000000000000000110110111000010001000000100111000001110000000000010000000000000011000001000000000000000010000000000001100000000000000000000110000000001110000100000000001010011000110100010000000000011000000000000000010000000010010000100000001000000000000001001100011000010011010000000011000100001101000000010010000000000100101001001010000100000000000000000000000010010000000000000000000000100111100010100000";
--X6Y9, LUT4AB
constant Tile_X6Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000100100001101001000000000100110011000011011001010011000000001110011000000100000000000100000010000000010001000000010000001001000000001100010000000110010011000000010001001100000100001100001111000000010000000000000001100001010000010000000000011010100001000000000000001000100000000011000001100001001001110110011000101100000000101001010010000110000101001000001000000011111000101001001100000010011001010011000001000000000100011000000000110000000100000000011001000000000001000000000001011101101100100001000110100001000100010110101000110000010000000001010001100111010001000000000111101001110011100100010000000000000100101000011010000100000";
--X7Y9, DSP_top
constant Tile_X7Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000011000000000000000000001100000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000001101000010100000000000000000000010111101101000000000000000000000000010100000000010010000000000000000110011110000000000000000000000000000001100000000000000000000";
--X8Y9, LUT4AB
constant Tile_X8Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000001000000001000101100000000001010101001000000111011111000001100011000010000001100000000000101000010000001111001011000000000110101100001100001110010000000001010000111010100101100001000000000110100001111010100000101101100000000000010100100000000000001111000000000000101000000000110101000000000001110000000000000100101010000000110000000000000101000001100000000000011000000100000100001010000010001101000110000101011000001000011110100100100000000101000100000000000100000001000001110000000001011111101011010000000010000000011110001000011000000000011001110100100101010001000000000100010111110001010110010000000000000100000000000000001110000";
--X9Y9, LUT4AB
constant Tile_X9Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000001000000001000000000000000110011001011011110000101000000101111011100000101000000010000010000010000000001001010100000001101100000000000001010000100100010010110001000010000000100101000000000010000000100000000000010000000100000000010000011000100000110000010000001100100000001000011010000000000000001000000000100000000000000100100000000100001001101000000000000000011100100000101011000000000000011100100000000010000000100000010101000000000000100000000000010000100100000100001000000000011010000101000000010001000000000110110100110000000000000000000100101100100000000000000000000000000111100011000000010000000000000000000000001000000000";
--X10Y9, RAM_IO
constant Tile_X10Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000001000100000000000000000000100100000000000000000000000000000100011000000100000000001000000000000000000011000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000010000000000000000000000000000000100000000000000000001000";
--X0Y10, W_IO
constant Tile_X0Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
--X1Y10, LUT4AB
constant Tile_X1Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001000101010000001100000000000000000000001000000000000110000000000001000000000100010000000000000100000000000000101000000100000000000100011110010000000110000001000001110000001000110000001000000000010001000110000110000010100000000010001100111000000000100000000001110100110000000000000000001000100011011101001000000100001000010110100000100111000000000001010000000000001000010000000010010000000010001011000000000000010000000000010000000000000000110000100000001000001000000001001100001101011000100100000001110000011100100010000010000000000000001000000001000000000000000000011100000101001010100000000000000000001000000000100011";
--X2Y10, LUT4AB
constant Tile_X2Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100010000100000000000010000001010000000000100000000001010001000010000000000010000000110000000000000100000011010000001000000011000110110010001010000000000010000001101100010100101001101000000000000000000010000111011010000010000000000001110000000000000000010000000000111000000000000000000000001110001011001110000000000000001010011100100001010010000000000000110011000000000110000000000010010000000000001010000000000000010000000100000001000000000000000000010000000000001000000000001000001100000011110100000000000110000110100000000010000000001010001000100011001000000010000110011000011001100010000000000000000000000000111000100000";
--X3Y10, RegFile
constant Tile_X3Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y10, LUT4AB
constant Tile_X4Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000111001000001000000000110011000111001000000000000001001110011100011110000000000000001010001001000000000000000000000000000000001000110000000000000000000000001100100100000000010100001000000000000100000001100001100011000000000001000000001001011001000000000000101000000000011100000000000000000000100001100110011000000000000010000000000000000010000000000000000101000000000000110000000001001000000000000000000000000000000000000000000000000000000100001000000000000001000000000010000000011111000010001000001000010000011000000000000010000000000010001010010000000000000000000000110000000000001110000000000000000000000000000000000001000";
--X5Y10, LUT4AB
constant Tile_X5Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000001000001000000000000100100010000000000111011111000001001010010000010001000000000000001010001000010100001111000000000000000100000000111110010101100010000000000101000000001100110001000000000000000000000000000010010000000000000011100100000101000000000000000011000000000000110100000000000000011000000010111000110000000000000000000010000000001110100100000000010000100000000001110000000000101011000000010000001000000000011001000011000000000000000000001001000000000000000010000000001000100110100000000010000000000000101010100100000000000000000001000100100100001000000000000001000110000000001000000000000000000000000000000000100010001";
--X6Y10, LUT4AB
constant Tile_X6Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100001000000000000101010000000111001100001000000001100010101100001111100000000000011010001001000110101111110000000001100100000000010010000000100010010010110000100100000000010100001000000001010000101010100000100001110000010100000100010000100111000000001000010100000100000110000000000000000001100000011000001000000000000011000010000100000100000001000000000000001000000001000000000010001000010010000000000010000000001110100000010000000010000000000010000000000000000000000010001101000101100000011000100000010000011000100000000000010000000010100011011000000001000000000001000000000000000000010000000000000000000000000000011000001";
--X7Y10, DSP_bot
constant Tile_X7Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X8Y10, LUT4AB
constant Tile_X8Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000100000000100000000001100000100000001000110000101001010000001101101011000001011111000000000010000011001000010100001001000000010100000111100000010010100000000110000100000101001100111100100001001100000101100100100000111101011000000000100000000000110100111000010001100010100010000000101000000000010000100110001111001101001000000000000000000000100001001011001000000100000000000000001111000100100001000001001000101000101000000000111000100000000000010000000000000011100000000100000000000000001100010101000011000001000010000100000100010000000010000000011010010101100010000000000000000000011011010011000010000000000000000000000001100101001000";
--X9Y10, LUT4AB
constant Tile_X9Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000111100001000000110011001001011011001011111000001100101001100010101000001000000010010000110010101000001000000000001100000000000110000011001000000010000000001000001000100100001000000000000000010000001000001011010010000000000100110011100010110000000000000000000100001011000000000000000001001000001100000000000000000100100000010000000001000000000000000001011110000000000000000100000000010000100000100000001000000001110000010100000000010000000000010000000000000000000100010000011010100110000011010100000000100000001100000000000000000000001111000000000111001000000000000010000010010101010000000000000000000000000000010011010000";
--X10Y10, RAM_IO
constant Tile_X10Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110100001111001000000000000000000000000000000000000000011100000000100000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000010";
--X0Y11, W_IO
constant Tile_X0Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000110000000000000000000000000010000000000000000000000000000011000001100000000000000000000000";
--X1Y11, LUT4AB
constant Tile_X1Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000001000000000001000100000000001010001001011001000000000000001100111000100010100001011010000011000000000010000000000000010001010001100001010000000000110011010000000010001000000000110000000000100100001000000100001011001000000000000010000000000000111001001000000000100001011001111110000000000000000000011000001110001111111000001010001000000000000001110010000000000001010111100000001111110000010010110001010000100010000000000000010010011110000001100000000000110011010000000000001000000001001010000111000011010000000000010010101000100000000010000100010101011000100010000100000000101110000001100000000000000000000000000100001011000000110010";
--X2Y11, LUT4AB
constant Tile_X2Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000010000000011110000000000000001010011000000100000000000010000000001000000000100000000000100000000000000000001101100000100000000011011010000000000010010100000000010001100001000000000000010001000000000100001010000010010100000000001100001000000000010001001000000011111000000000001100000100100010000101000000000001000000000100100000001000000000000000000000000000000110000000000000000000001100001000000000000000000000000100100000000000000000000000000000001000010000000000000000001100000000100100000010000000000000100110000010000000001010011000000011001000000000000100100001011001000010000000000000000000000000000000000010";
--X3Y11, RegFile
constant Tile_X3Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y11, LUT4AB
constant Tile_X4Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001000000000000101011111000000000101000010000000001010000000010001011000000100000010000010010000100001011010000100000100000000110010000010000000000000010001000001101010101101001000000101000110010001001000110001000000010111101100000101000000000000001101101000000001010011010000000000101000100000011010010000001001001011000010000001100011100001101000001001001000000100011000000010100000010011000100111000100000000101000000000000001100010000001000000010000000000001000000001000100010100000000010000000011100100000100100000000010000000000000001000100001000000000000000000000010000111100000000000000000000000000000000010000000";
--X5Y11, LUT4AB
constant Tile_X5Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000011111000000110010101001111000000000000000001100100010010111100000000000100001110011100001001100000000000000000000100000110110000000111000000000000100100000000001100101001000000000001101110000000010001010000000000000111000000000011000000000000000011101010000000010111000000000000110010010001010000000000000000000000000000101000000101000000000000001000100100000001111000000000100001000010010000000000001100010000000000000000000100000100000000000000000000000000010000000000010000000010000100000000011000001101101000100010000000000011111001001111000001100000000001100110001000000100010000000000000000000000000000110000000";
--X6Y11, LUT4AB
constant Tile_X6Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000101000000100000000000000001000100000010111110001100000000000010100000100010101001000000000010010000000010100100011010000011100000011110000100001111000001010000110000010000000100011100001001100101111010101001000000100001000000010101100100000100001110000000000011000000000001000000000000000001110000100000000000000100000000000011000000010110001100001000000000000101000010100001001100000010100010001010010001000000000100011110100001100000000100000100000100011000001001000000010000000010000001010000011010000000010010010101000100100010000000000011001110000100000000000000000100000111001000000000000000000000000100100000000100011010001";
--X7Y11, DSP_top
constant Tile_X7Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010100000111010100000000000000000000000000000000010010000110100000000000000000000000000000000000000000000000000000000000000000000";
--X8Y11, LUT4AB
constant Tile_X8Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000001000100000000000011111111000100100000000000000000000010000110001111100010010000100010000001000000001111000000001010000000011100100000111000000011100011000011010000000001010000000101110100000100000100000101000000100000100011000010000000000000000010000010001010000100101001000000000000010001001001100110000110000000110001000010001001000001001000001101010011001001000100111110000000001110100000000000010001000110001100111010101001000101000000001100100100000000000001100000000001001100011100000000001000001010010000000000000000000000000011101100000000001000100000000000010000110011000110010000000000000000000001000001101000010";
--X9Y11, LUT4AB
constant Tile_X9Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000101000000000000000010110000000000000001000010000001100000001000100001111001000000001110011000100000001111110010000000000100000100101110000101000000000100001101100001000100101001000000000110000110100001000001010000100000000000100100011000001001000110000001000101000000001011000010000001001000000001000000101000100010000001010000011101000111000001000101000000101000000001010000000000110001100000000101000011000010011100101001010000001000000000000000010010000000000000000010001010000011101000000000001000011000101101100010000010000100000001001000001000111100000000000001000001001101000000000100000000000000001000011000100111000";
--X10Y11, RAM_IO
constant Tile_X10Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001010000010110000000000000000000001101100111100000000000000000000000000000000000000000000110000000000100000000010110000110000100000000000000000000000000011100101111101010000000000000000001010001000100010101100101010110000001010000000001000000011111101010100100000001010001111001000";
--X0Y12, W_IO
constant Tile_X0Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000011100001110000000000000000000000";
--X1Y12, LUT4AB
constant Tile_X1Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000110011000000110100000000000000010011010000001100000010000000000011000000000101100001100000100100000110000000100000000000000010000010011010000000000010100001000000000101001000000010000010010000000000001011010100000000000100000000001010110000010000000010000000000011111000000000000001000000000011010100000000001100000000011110010000001000001000000001000000000000000111010000000000000110110000010000100000000011010010011110000000010000000000010000100000001000010000010000000100000001000011000100000000000110100101100110000000000000011000011011010110001000000000000100000101000000100000000000000000000000100000001001010000";
--X2Y12, LUT4AB
constant Tile_X2Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001000000100000000000001000001010000000000000000000100000000000000100000000000101100000000110110000100010000001110001000001101000000000000100011000000000001100100001000110001000100100100000110001000101001010000000000000000100110001111000110000011000101100011010000001100000000000101001001010000011111000100010000000101000001111010100100101010000000001000101000001001001111000000100000010010000100101001000000010010100010001110000100000100000101000100000010100000000000000010100000010010000110000000001010010101111100110000000000000011101010011010101001100000000000100000101010001100010100000000000000000001000001011000000";
--X3Y12, RegFile
constant Tile_X3Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000111000001110010000000000000000011000000000000000000000000000000";
--X4Y12, LUT4AB
constant Tile_X4Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000101001001100000000100001111001000000000001111000001000110101010011110111010010000001010101001011111100100111000000100001100100010010100011001000000110000000100010100000011100101001000010000000000110011100011011011100000000010000000000001010000000000000010001000000001011000000000000000010000110101111110110001000000100000010000000000001010001000000000000000000000010000110010000000010000011100000000000000000000011010000000100001001000000000000100100100000000000010000000001010100000000000011010000000000010000000000110000010000000000000000000110000010000100000000011010000100000001001000000000000000100000001000100011010000";
--X5Y12, LUT4AB
constant Tile_X5Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000111000000001000000000000000000111000010000101000000000000000000001100100010010000001010111000000110100100001000000000000000111100110000000001000000000000011111100001100000000100001000000000100110000010100001100001100000000110000100100010001001000000000000000001010111001110000000000000101000100000000001101010000101010000000010000001001000000000000000001001000100000100000010000000100100000000010000110000000110011100000000000000000000000000000000000000000000000011000000000000000000100000000000100000011000110001100100000010000000000010100001100000000000100000001001000010000000001000000100000000000000000000001000000010000";
--X6Y12, LUT4AB
constant Tile_X6Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000001000000100010000000000000100000000000000000010010101000000001100001000111100101010010000001100000010000101000100011000000010001100011100010100011000011000000000110110111100000010010000000001110001000100100101100011001010100000010101001110001001000000000000000101101000000001110000000000000010000000010101011000110100000001100010100000000010001010111000000000000000000100000100111100100000011000010000000000001000001000000111000000000000000100000000000010000100000100000000010000000100100000000000000000001000010011011010100100000000000000010000000011111000010000000000000000100000100000000000000000000000000100000000000100100011000";
--X7Y12, DSP_bot
constant Tile_X7Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010100000000011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000";
--X8Y12, LUT4AB
constant Tile_X8Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011010000000111001000001111000000100001001000001110001010000100001000011000001001100100010000000010001000010000000100001100010010100000111010001000001111010001001100100101000010100001011000010001100000010110100100001111000000000100001101001000000100010000010000000110101010000101000011000011000000010100000011111001000000000001001001101000010000000101111010000000100101100110000000010000100010000000000000100000000101000000000000010000000000000001000000000001000001000000111110000000001000111000011100000010000100000001110000100010001001100000000000000000010000000000000000000000000000001000000000110011000";
--X9Y12, LUT4AB
constant Tile_X9Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000010001000000100000000000000000000000000000000000000000000000000000001010000000000000000000000010010000001001000000000000000000000000010000000000000000000000001000001100000000000000100000100000000000000000000000000000000000000000000000000010000000011100000000000000000000000000010000100000000000000000010000000000110100000000000000000000000000100000011000000000000100000110000000000000000001000010000000000000000001000000000000000000000000000000000100000000000000000000000000000000011010000000000001000000000100000100000000010000000000010000000010100100000000000000000010000000000000000000100000000000000000000000000000001000";
--X10Y12, RAM_IO
constant Tile_X10Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000110010010001000000000000000000000000000000000000000011000000010000000000000000000100000000110000000000000000000000000000000000000000000000000000000001010111111101110000000000000000001010001001011000011111011010100000000000000011000000001111111100000000001010111100101011001010";
--X0Y13, W_IO
constant Tile_X0Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000011100011110111000000000000000000";
--X1Y13, LUT4AB
constant Tile_X1Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000001000000000001000000000000000000000000010000001000000000000000000000000000100000010000";
--X2Y13, LUT4AB
constant Tile_X2Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000";
--X3Y13, RegFile
constant Tile_X3Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y13, LUT4AB
constant Tile_X4Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X5Y13, LUT4AB
constant Tile_X5Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000";
--X6Y13, LUT4AB
constant Tile_X6Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000010000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000";
--X7Y13, DSP_top
constant Tile_X7Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X8Y13, LUT4AB
constant Tile_X8Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010010000";
--X9Y13, LUT4AB
constant Tile_X9Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010100000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X10Y13, RAM_IO
constant Tile_X10Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000010110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000011000000";
--X0Y14, W_IO
constant Tile_X0Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101101110100000000000000000000";
--X1Y14, LUT4AB
constant Tile_X1Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001110000000000000000000000000000000000000000000000000000";
--X2Y14, LUT4AB
constant Tile_X2Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X3Y14, RegFile
constant Tile_X3Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y14, LUT4AB
constant Tile_X4Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X5Y14, LUT4AB
constant Tile_X5Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X6Y14, LUT4AB
constant Tile_X6Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y14, DSP_bot
constant Tile_X7Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X8Y14, LUT4AB
constant Tile_X8Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X9Y14, LUT4AB
constant Tile_X9Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X10Y14, RAM_IO
constant Tile_X10Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011";
--X0Y15, W_IO
constant Tile_X0Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000011100001111110000000000000000000";
--X1Y15, LUT4AB
constant Tile_X1Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000110000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000";
--X2Y15, LUT4AB
constant Tile_X2Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X3Y15, RegFile
constant Tile_X3Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y15, LUT4AB
constant Tile_X4Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000";
--X5Y15, LUT4AB
constant Tile_X5Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X6Y15, LUT4AB
constant Tile_X6Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y15, DSP_top
constant Tile_X7Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X8Y15, LUT4AB
constant Tile_X8Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X9Y15, LUT4AB
constant Tile_X9Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X10Y15, RAM_IO
constant Tile_X10Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y16, W_IO
constant Tile_X0Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101111110101000000000000000000";
--X1Y16, LUT4AB
constant Tile_X1Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000";
--X2Y16, LUT4AB
constant Tile_X2Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X3Y16, RegFile
constant Tile_X3Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y16, LUT4AB
constant Tile_X4Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X5Y16, LUT4AB
constant Tile_X5Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X6Y16, LUT4AB
constant Tile_X6Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y16, DSP_bot
constant Tile_X7Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X8Y16, LUT4AB
constant Tile_X8Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X9Y16, LUT4AB
constant Tile_X9Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X10Y16, RAM_IO
constant Tile_X10Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
end package emulate_bitstream;