// X0Y1, W_IO
`define Tile_X0Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y1, LUT4AB
`define Tile_X1Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X2Y1, LUT4AB
`define Tile_X2Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X3Y1, RegFile
`define Tile_X3Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y1, LUT4AB
`define Tile_X4Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X5Y1, LUT4AB
`define Tile_X5Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X6Y1, LUT4AB
`define Tile_X6Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X7Y1, DSP_top
`define Tile_X7Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y1, LUT4AB
`define Tile_X8Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y1, LUT4AB
`define Tile_X9Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y1, RAM_IO
`define Tile_X10Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y2, W_IO
`define Tile_X0Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y2, LUT4AB
`define Tile_X1Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X2Y2, LUT4AB
`define Tile_X2Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X3Y2, RegFile
`define Tile_X3Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y2, LUT4AB
`define Tile_X4Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X5Y2, LUT4AB
`define Tile_X5Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X6Y2, LUT4AB
`define Tile_X6Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X7Y2, DSP_bot
`define Tile_X7Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y2, LUT4AB
`define Tile_X8Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y2, LUT4AB
`define Tile_X9Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y2, RAM_IO
`define Tile_X10Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y3, W_IO
`define Tile_X0Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y3, LUT4AB
`define Tile_X1Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X2Y3, LUT4AB
`define Tile_X2Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X3Y3, RegFile
`define Tile_X3Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y3, LUT4AB
`define Tile_X4Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X5Y3, LUT4AB
`define Tile_X5Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X6Y3, LUT4AB
`define Tile_X6Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X7Y3, DSP_top
`define Tile_X7Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y3, LUT4AB
`define Tile_X8Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y3, LUT4AB
`define Tile_X9Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y3, RAM_IO
`define Tile_X10Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y4, W_IO
`define Tile_X0Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y4, LUT4AB
`define Tile_X1Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X2Y4, LUT4AB
`define Tile_X2Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X3Y4, RegFile
`define Tile_X3Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y4, LUT4AB
`define Tile_X4Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X5Y4, LUT4AB
`define Tile_X5Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X6Y4, LUT4AB
`define Tile_X6Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X7Y4, DSP_bot
`define Tile_X7Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y4, LUT4AB
`define Tile_X8Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y4, LUT4AB
`define Tile_X9Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y4, RAM_IO
`define Tile_X10Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y5, W_IO
`define Tile_X0Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000011000001100000000000000000000000
// X1Y5, LUT4AB
`define Tile_X1Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X2Y5, LUT4AB
`define Tile_X2Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000111110000010100110000000000000000000010000000001100000100000000011000000000010000000010010000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000001010000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000011000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000
// X3Y5, RegFile
`define Tile_X3Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y5, LUT4AB
`define Tile_X4Y5_Emulate_Bitstream 640'b0000000000011000000100000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000100000110000000000000000000000001110000000000000000000000000000000000000000000000010000000000000100000100000000000000110000000000100000000000000000000000000000000000000001000000001100000000010000000000000000000000000000000001000000000000000000000000000000000000000000000001010000000000010000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000
// X5Y5, LUT4AB
`define Tile_X5Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000100000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X6Y5, LUT4AB
`define Tile_X6Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X7Y5, DSP_top
`define Tile_X7Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y5, LUT4AB
`define Tile_X8Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000
// X9Y5, LUT4AB
`define Tile_X9Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y5, RAM_IO
`define Tile_X10Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y6, W_IO
`define Tile_X0Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000011101001111111000000000000000000
// X1Y6, LUT4AB
`define Tile_X1Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000011000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000
// X2Y6, LUT4AB
`define Tile_X2Y6_Emulate_Bitstream 640'b0000000000000000010100000000000000000001000001001001000010001000000100000000100000000101000000100010000000000000001100000000000001001001100000000100000000000000011000100100001000100001001100100001110000001001010100001100100101011000000000000000000001101111001000101001100001000000001011001000000000000000001000001111000001100000000100001000000000100101001101000000000001010010100000000110100000000000011000000000001101000000000001100000100000000000000000000000000001100000000000000000000001001000100100001000000000000000100010000000100000010010000000000010111010000001000100000000000010111100011010000000000000000000000000000001000100000000
// X3Y6, RegFile
`define Tile_X3Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000101001000000000000100001001100000000001100000001010100000000010000000000111000001001001010001011110010001110001100001100001011100000000000001100000000000000000000111010000000000100000001000000010000000000001100000000000000100000000000100000010101011111000010011011000000001101100010100000101000000000011100000100000000000000000011000000000000000000000000000000
// X4Y6, LUT4AB
`define Tile_X4Y6_Emulate_Bitstream 640'b0000000000000001111001000000110000010000000001110011000000000000000000001111100001110111010010000000010111101110101000111110000000000100000100000010100001001000000001000010001110000001010100101001100100000110010101101101000110001100000000100000110100100000000001010000000001000000000001010000001100000100000100010000000010000001000000101000011111001000000000011100000001100100000000000000001000000101011000000000000000101000000001101000101001000000001000100000000000000000000000000010000000001010011001001000110000000011100000000101000010000000000000000000000010110000000000000000000100101000000000001010100000000000000000001001000001100010
// X5Y6, LUT4AB
`define Tile_X5Y6_Emulate_Bitstream 640'b0000000000000000100000000000000000000001010001000110011010111000000101000010010000000000001000100001100010000000010001100010010000011100100011101001100010000000000010000100101000000100100110000000000000101101000000001000010000000110000010100000100001001000110000100001101000000000000000000000000000000010001100001100000110001100000000000000010000100100010100000000000000110000000000000000000000010100010010010000001101000000000011010000011100000000000000000000011000000000000000000000000001101001000000000010000000000001000101101100000000000010000000010010011101100100000100000000000000111000100110000000000000000001100000001001000000000000
// X6Y6, LUT4AB
`define Tile_X6Y6_Emulate_Bitstream 640'b0000000000000000111000000000000000000000000000100000001001010000000001100001010100010000001000000000000010011000000000000000000000001000000011100100000000110010000001010000001000100000100011100001001001100000100001001000000100001000001000011000000001001000000000000000001100000001000000010000000000000100010000011100000000001000000000100000000000001001100000000000000010000000001000101000000000000101000000000000000010000000000000000000011110000001000000100001000000000000011000001000000001001010000011000010000100000000000000000000100100000000000000010000000001000011000100000000000000000000000000000000010000000000000000000000000000010000
// X7Y6, DSP_bot
`define Tile_X7Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001110000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000010000000000000000000000000000000000000000000000001000100110001000100010000000100000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y6, LUT4AB
`define Tile_X8Y6_Emulate_Bitstream 640'b0000000000000000000001000011000000001100110000000000010010000000000001100011000010000000101110000000000000000010110100000000010000000100100000001010000000000000000000010000000010000000000011000000000010000000110000001001111000000100000000001100000001101001001000000000000101110000000010100000000000010001010000000001110011000000000100001000000010100100010100000010000100000001000000000110000000000100000000100000101101001000000000000000101001000000000100100001000011100010000000000100000001000010111010000010010000000001001000000000100010010010000000001000000001000100000000000000001000000111001001000010000000000000000000001000000000010000
// X9Y6, LUT4AB
`define Tile_X9Y6_Emulate_Bitstream 640'b0000000000000000011000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000010100100000000000000000100000000000010000000000010000010000000001000001100000000000000000000000000110000000100001000000100000000001100000000001000110000000000000100011000000011000010000000000001010000000011000100000000000000011000000000000000000000000000000000000000000000000110000000000111010000000000000000000000000001000000000000000000010000000001010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001000010000100000000000000000001010000000000011100000100000000000000000000000010000000000
// X10Y6, RAM_IO
`define Tile_X10Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000100000000000000000000000000000001100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000
// X0Y7, W_IO
`define Tile_X0Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101011110100000000000000000000
// X1Y7, LUT4AB
`define Tile_X1Y7_Emulate_Bitstream 640'b0000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001001000000000000
// X2Y7, LUT4AB
`define Tile_X2Y7_Emulate_Bitstream 640'b0000000000000000000000010101000000010001000000101000000001111000000000000000010000100010000000000001100000110000001000000101000000000101000000100100100000101011000010000100100000000001100101101001000000100001000100000001000110001000000010010000000000100000110000011000010000100010001010111000000000000000000001000000000000110000010100001000011111110001101010010000000010000001000001001000101000010000011010000000101100101010000000011101101000000000110000000000010001110000001000010000010000010110111100011000010100000001000010110111100000010000000000001001111110010100011000000000001100001001001001000000000000000000100000001000000011110000
// X3Y7, RegFile
`define Tile_X3Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000110010011010000011000000000100010000000000000000000000000000000000011011000100000000000000000000110110100001110001000101111000010000100111000000100011000000000000111000000000001001001100010010000000000000000000000000010000001001000000000000000000000010001000100000101100100001000000111001100001110111010000010000000011110101000001110111100000000000000011000000001100000000000000100000
// X4Y7, LUT4AB
`define Tile_X4Y7_Emulate_Bitstream 640'b0000000000000000000101000000000000000000000001000000110000000000000001101101010110000000110100000000000110000001011000000000000000000000000101101010000000100000000000100000001000100100100000000000000000100000110000001100010000000000000000001100000001000000000000010000000000100001001000000011000000000000000000001000000000000000000010100000000011100001100000010001000000000000100000001110001000000000100000000000001000000000010001001000100100000001000000000000001011000000001000000100000001100110111000011000000000000010100100000000000000010000000000000000000101000000000000000000000001110000000011010010000000000000000000100111100100110000
// X5Y7, LUT4AB
`define Tile_X5Y7_Emulate_Bitstream 640'b0000000000000000000001110000000000011111100001011011111010000000000000000011000011100101101000000001000000000011001000000111000001000000000011000101100000000000010000000111101000000000001100000000100010001010110100001010010100000000000010110101000100010010000000000000001100000000000001000010000000010001001001010011010000000000000000000000010000101000000010000000000001010110100000100110000000010000000010010000001010000000000000101100001000000000000000100000000110000000001100011000000000000100001110001000100100000001000110101101110010010000000000011110001100101101001100000000000101101000000001000000100000000001000000000010001100000000
// X6Y7, LUT4AB
`define Tile_X6Y7_Emulate_Bitstream 640'b0000001000000000000001110000010000101010000000000000101000110000001000101000100001100100101010000001010000000000100000100000010000000000000001011110100000000011000001000100001000000000010000000000000100001001000101101000001101010100000010001001010001110010000000000000100000000101011001000010000000010100010000100011111000100000001000101000000011110000000001000000000000000101000000000000100000010101000010101000100010010000000001001010000000000000000000100001001010000000001000001000000000000000000000010000010000000000110110000110100010000000000000000010001011101011000000000000000000000000010001110000000000000000001000001010000101000000
// X7Y7, DSP_top
`define Tile_X7Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000110100000000000000000110010000000000000000000000001100000000000000000000000000000000000000100000000000000000000000000000000000001011000000000000000000000000000000000000000010100000001011100000000010100000111100000000101000000000110011010000000000000000000000000000000000000000000000000000
// X8Y7, LUT4AB
`define Tile_X8Y7_Emulate_Bitstream 640'b0000000000000000100000000000000000000000000000000000100001100000000001100010100110000000100100100100000110110000000000100000000000101000000000100100000000111000000010000100010001101000111000000000000010100001000010010100101000000110000000000001001000011100110001001000000000001100011010011010000000011100011001000000000100000000000000011010000000010001001011001000000010010111110000000110000000000000000010000110010000000100000000000000000010000000100000000000010000000000100000010000000000001000000000000001000000000000000010000000100000000000100000011000001100000001000000000000000000000001100000100000000000000000000001000000000000010000
// X9Y7, LUT4AB
`define Tile_X9Y7_Emulate_Bitstream 640'b0000000000100000010000000000000000010101010000000000000000000000000000001000000100000010100100100100000000000100000000001000000000000000000111100010000000000000010000000110000100001100000111000000110000100011000000101000000100000100000000001100000011000000000010000000000010000000100001011000000000010001000000000110100000000000001100000010000000000000001000001000000100000010000000000000000000001001001000000000001100000010000000000000000001100000000100000001010000010000000000010000000001000011000001000010000100000011000000011100000000010000100000001011000000000010000100000000110000100010100101110000000000000000000001000111011000000001
// X10Y7, RAM_IO
`define Tile_X10Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000001111000000000000000000011000000010000000001010000100000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010
// X0Y8, W_IO
`define Tile_X0Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110110000000000000000000
// X1Y8, LUT4AB
`define Tile_X1Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000100000001000000000000000000000010000000100000000000000000000000000000100000000000000000000000000000000010110000100000000000000000000110000000001100000000000000000000000000000000000000000
// X2Y8, LUT4AB
`define Tile_X2Y8_Emulate_Bitstream 640'b0000000000000000000001010111100000000001010000100100010010111000000001000000010010010001010010000001110000010100010000000000010001000000000011100010000001000011010100000001010110101101000011001001111000001001000000000101011011011100000010000000000000000011001010110001101101100000100001111011100000000010001100000000011011101001100111000000010000000100011010001100010100010000100000000110110100010000111111111000000000010100000000010100000010000000001010100001100000110000001100010001000001101100010100100000000111000000101111001111100000000000000000001001010000010011001000000000000100000101010100001010000000000000000000111010000001101000
// X3Y8, RegFile
`define Tile_X3Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000101000000000110010000100000100100000100101100000000000000000000000000000011100010011011000000000000000000000010000010111000000000001110010011011000011110111000010000100110000000100000000000001000100011100000000000000000001000000010000001000000010000101110100100000000010110010101000100101000000000001100010001000011101010001000000000000000000110110011100100000000011000011001100000000000000100000
// X4Y8, LUT4AB
`define Tile_X4Y8_Emulate_Bitstream 640'b0000000000000000101000110000000000001010000001000111010010011000001100001101010000010111010000000001100010001001111100100111010000011001100000000010000111000101000000110001100010000000010000000000101100000000010001100001001001010000110000000100100010000001001000000001101100000001101000100000000000011100000000011100000001001100000100001010000001110001100011100010000101000001000001001001001000000110000010010000001100001000000000110100111100000000100000000000100000000000000100010000000001000101111110000000100000000000000000001111100011000000000000010101001001001000000000000000000011110111100010000000100000000000100000010011001000000001
// X5Y8, LUT4AB
`define Tile_X5Y8_Emulate_Bitstream 640'b0000000001000000000010000000000000100000000000010000101000000000001100100101000000100011101000000110110001000000100000101011000000000001100000111110100000000011000000010011011000001100000001000000101000100010010000000101001000000001000000000100100000000101001000100000000111000010100110011000000010001101010000101100110101100001001000101000000011010001001101000110011001000001101001000001100000000000000000010001000001101000000001110000001010100000110100100001000000100000001000010100000000000010111111000011100100000001100111010101100100000000000000001110000010001010001000000000001110000001001010100000100000000000000000001000000011110000
// X6Y8, LUT4AB
`define Tile_X6Y8_Emulate_Bitstream 640'b0000000000000000010011110000000000011001100001111000101010000000000000000000000001110011000000000000000000001000101000010111000000001101000010000010010001000010011010100101110100100000001000000000001000001001110100000100010001010110000010000000100111000100111000000001101110000000000100000001000000000010001000110011000101100000001000101000010011110000000111000000000001010001000001000000100000010111001110010000000001001000100010010011000100000000000000100000101100000000000000000100000001001110001111000000000100000011000010110100000010000010000000011001000011101100010000000000000000000000110100000000110000000000000000001001001001110000
// X7Y8, DSP_bot
`define Tile_X7Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000110000000000000000000000010000000110011001100100011000001100011000000000000011000000000001000000000000000000000000000000000000000000000000000000000000000000000
// X8Y8, LUT4AB
`define Tile_X8Y8_Emulate_Bitstream 640'b0000000010001000000000000011000000010001100001111011000000000000001100001000000101011001001010100000000010001110000001011010000000001000000000010000100001000011000100010010001010100000001000000001110000100110110100001100000100001000000000100000000111010000000010000000000000001110001000100010100000001100000100010000100100111000000101000010011100001000000010000000000000000001000000100000100000000001000000010000010010001000000000010101000110000001000000000000000000100000000000001000000001001000100001001110100000000000100010001111110000000000000000000101100011101000011000000000000000000100000101100010010000000000000000010010001000010000
// X9Y8, LUT4AB
`define Tile_X9Y8_Emulate_Bitstream 640'b0000000000000000110001001110110000000000001000100100010000100000000000000000110010111110000000000000000001000010101100001010000000001101000110000110010000010100000000010100101000000000111001000000110000000100000100000001000000010000000000110001110100111010000000000000101010100010000011111000000000010100100000000011010010000000001100100000000001001001110000000000000000000011000000001110000000000101010010000000000000001000000001000000000001100001000000000000011000000000001000000100000000010000100010001000110000000000000000001111100100010000010000000101110000100100001100000000011100100100000011101000010000000000000000010000000000001001
// X10Y8, RAM_IO
`define Tile_X10Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000100011110000000000000101011000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010
// X0Y9, W_IO
`define Tile_X0Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000111100101110000000000000000000000
// X1Y9, LUT4AB
`define Tile_X1Y9_Emulate_Bitstream 640'b0000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000011000000000000000000000000110001000000001000000001000000000000100000000000101000101100000000000000000000000010000000000000000000000000000000000000000000000000000011100100000000000000000000000010000000110000000000000000000001000000000000000000000000000000000000000000000000000000000
// X2Y9, LUT4AB
`define Tile_X2Y9_Emulate_Bitstream 640'b0000000110000000110000110000000000000000101001110000000000000000001100101000010100000011000000100011000001000100000100000000000000000001100100010000010000010000010000010000100101000000010000000000000000000000000100000001011000000000000000010001000000100000000000011000010011100000010000000000000000001010110010001101001010010010001001000000000010110100000101000001000110000100000001000000000000000001001010110000101111000001100010001101010000000001100100000000000000100000000000001000000001001010001010000011010000000010000100000000110010000000100000000111011100001100110100000000000010100000001000010001010000000000000001010001000110000001
// X3Y9, RegFile
`define Tile_X3Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101010011011000000000000001010100011100000000000000000000000000000010011011000000000000000000000111010001001110101000101111001010010001100001000000011000100000011000000011000100101000000000100000000000000000000000000000000010000001100001001101000001011000001110001110110000000000011100011001001000111011100000000001000000101010000100110010100000000000011000000000000000000000000110000
// X4Y9, LUT4AB
`define Tile_X4Y9_Emulate_Bitstream 640'b0000000000011000011110110100000000000110000000100100000001010000000000000011000101011101000000000010000001001100000100001011000000000001000000000000100100010110000010010000100101101100100000000000111000000011010100000100001000000100000000000100001000001010000000010000000011000000100010100001000000000000010010101111000000000000000100010010001110100000000001001101000000001100001000001111000000010000011001000000111100000000000000100000000100000000100010000000100001100000000100010000010000001010000001001000000001000010010100000111000000000000000000000010111000100000011000000000000011001111010100100010100000000000000000011000101110000010
// X5Y9, LUT4AB
`define Tile_X5Y9_Emulate_Bitstream 640'b0000000000000010001001110100000000100000000001111000000001010000000100000000110000101011000100000110110000000000101000001011010000100001100011101110010000000011000000010100011000001100000010000000100000101001000000000000011100000000000000000000110010110000110000010000001001010010100101000010000000001100010100001010100110101000000001001000001101000001010100001000000010001001000000000000100000000101001100110000001001000010000001110011000110000000010000100100000000100000001100000001000001000000000101010011010010000001000000100111000100000000000100011111111110101000000000000011000010000011001000000010000000000000000000000001100000000000
// X6Y9, LUT4AB
`define Tile_X6Y9_Emulate_Bitstream 640'b0000000000000000000001100010000000000110000001010011111011100000000100000101100111100001101100100111010000000000011100000000000000110000000011101110000001010010010000000000111001000000101010000000010001100000110000110001000000000100001010010000010100100000110000000001101100000000100000000000000000000101010000100011010100000000000000010000011100110100000000000000000000000100000000000001010010010100001010010000110000000001000001010001000100000000100000000000110000100000000000010000100001010110001100100111110100000011000000100110000000000010000000010011000010100000001100000000000000000000100011000000000000000000000000000000000000000000
// X7Y9, DSP_top
`define Tile_X7Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100100000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000001000000000000000110000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000101000001011000000001010111000000000000000000000000000001110110000000000000000000000000011110000000000001010000000000000000000000000000000000011
// X8Y9, LUT4AB
`define Tile_X8Y9_Emulate_Bitstream 640'b0000000110000000100000100000000000000000011000000000001010110000000100000000000010001010001000100101000010000000010101011000010000100000100000101010000001110101000000000000101010100000010010000000100000000111000001010100010000000010000000000001010100000010110000010000100001000000111000110001000000010000010000011000000110000010001000000010011000110001110010000000000011000000000101101001010000010001000000100000011000001000000001010100110000000000100000000000010000000100100101000000000001010011100000000001000000000000000010100100000011010000000000000011001001000100010000000000011101110010001011110010000000000001000000000000000010000000
// X9Y9, LUT4AB
`define Tile_X9Y9_Emulate_Bitstream 640'b0000000000000000001000000000000000000000000001000010010000100000000000000000000000000000000000000000010000000010110100000000000000001100000000001010000000000000000110100010001000100000000000000000000000000010000000000100000000000100000010000000000010100000100000000000100000000001110001000000000000010000000000000000100000000000000000000000000100110100000100101000000000000000000000000110000000010000011010000000001101000101000001000000000100001000000000000000000000000000000000000000000000010011011000000000010000000010000100000000000010000000000000010100001000000000000000000011000000010000000000000000000000000000000000000110000000000000
// X10Y9, RAM_IO
`define Tile_X10Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001111000000000000000001100000000000000000000101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000
// X0Y10, W_IO
`define Tile_X0Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010
// X1Y10, LUT4AB
`define Tile_X1Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000001000000011001000000000000000000000000000000110000000000000000000000100010000000000000000000000001100000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000100000000
// X2Y10, LUT4AB
`define Tile_X2Y10_Emulate_Bitstream 640'b0000000000000000011000100000000000000111100001010011001010000000000000000011100000100000001000000001010000010001001000000000000000011001100000010000000101110010000000000000100000000000110011000000001100000100000001000000000001010010000000101101010010000000000000010000000000010010000011000010000000000001101000100011010010001000000000000000000000111100110110001001000100001010000001101010000000000010000110111000001111000100010000001010010110000001100000100001010111100011001100001000000001010010100001001000000000000000100111100100000000000010000000000100111010000010000000000000001100000000001010000000000000000000100000000011000110000010
// X3Y10, RegFile
`define Tile_X3Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000110010101011000011110000100000000010010000000000000000000000000101100101001000000010000000000000110000100001111000000001101100010100110000111111111100000000110000101100000100000000000001110000000000000100000000000000000000111000011100000000010110101010000010001000010101010111110000001101100001100000011000010000100000000000000000110010000010010100011000000000001100000000000000000000
// X4Y10, LUT4AB
`define Tile_X4Y10_Emulate_Bitstream 640'b0000000000001010111100000000000000011110000001100010100011001000001101100000000001010000001000100011010001011000111100001000010000010100100010010010000001000110010010100000011111001000011010000000000100000000010000010000011000000100100000000000010000110000110000100101100010111010100001100000000000000000000000110100010010010100001101001000000111011000010000100101000000101111100001001001000000001010000001010000101000000000000000110001100010000000101000100000110011000000000100000110000000001010011000000100010000000010110001100100000010000000000000010000010001000000010000000000000000000101001011000000000000000000100000101001101000001000
// X5Y10, LUT4AB
`define Tile_X5Y10_Emulate_Bitstream 640'b0000000000000000110101100100100000000001100001111000001010000000001000000000110001100010010000000001000000011000010100011100000000001000000000010000000001000110001110000010000000100000000000000000100000101000110010001100000000000010000010100001000001000000000000010001100000101011101011110000000000001100001101010011000000100000001000001000011101000101000001000001000010010000000001001000100001010000011010000000000000000000110000001000000100001001010000000000100000100000000000010000010000101110000001100011000000000001010010000111100000000000000000010101100011000000000000001000001011110010110000010000000000000001000000000001100010011000
// X6Y10, LUT4AB
`define Tile_X6Y10_Emulate_Bitstream 640'b0000000000000000100111111000000000001010101000000011001010011000000000000000000100001010010110100000010100000100000000101010010000001101000110000110110001010010010000000010011110000000001011100000000000000110100000001001010001010110000010110001100000010110001000010001101100000110000101000000000000000001001001100011000011000000001000000010000100011000010011000000000000000111100010100001000000010000000011011000101110001001000001000100001100101000100000000011000010000011000000011000001000000101110000101001100100000010000000100000001010000010000010011101001010000000001000000010001000000001111001111010010000000000000000010000100110000000
// X7Y10, DSP_bot
`define Tile_X7Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000110001001100000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000110000000000000000000000000000000000000000000000000000001000000000000001100000011101110000000000000011000000000000011101000000001000000000011100000000000000000010000000000000000000000000000000000000
// X8Y10, LUT4AB
`define Tile_X8Y10_Emulate_Bitstream 640'b0000000000100000100011000111000000000000000000000000011010000000001100001000000000000000010000000011000110000000000000001000000000101001100000000000000101001000010000000000100001100000000110000000000010100101100011110100000010000110000010011101001000000000000000000001110000110000000000110010000000011000101011000000111100000100000100000010010000111000010011000000000110010001000001000000010000010011010110101000111000110000000000110001000010000000110000000000001100000000000000000000010001010011000001001000000000000000011000000000100000000010000000001000000000000000000000000000101001110111011000010000000000000000100100110001100000101000
// X9Y10, LUT4AB
`define Tile_X9Y10_Emulate_Bitstream 640'b0000000000100100010100000100000000010100101000110000010010000000000000101010000101100000000000000000010110100100000000000000000000010100000101110110000000000011000010000010011100100000000100000000000000000010000000000010000001010000000010000001000001000010100000000001000010000000010001000001000000000000100000001100001000100000001000000010001011010001000000100001100100000010000001000000100000010010010000001000000110000100110001000000000100010001001000000000000000000000010010001000000000000011000000000101100000000011000100000000010000010000000000000011010110011011011000000000100000000000010000100011000000000000000000000001100000101000
// X10Y10, RAM_IO
`define Tile_X10Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000001000000000000101000011111111100000000000000000000000000000000000000001000001100000000001000001000111100000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101010101000001000100000000000
// X0Y11, W_IO
`define Tile_X0Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000011000001100000000000000000000000
// X1Y11, LUT4AB
`define Tile_X1Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000010000000000000100000000000110011000000000001100000000000000000000000000000000000000000000000000000000000000
// X2Y11, LUT4AB
`define Tile_X2Y11_Emulate_Bitstream 640'b0000000000000000011101000000000000001010101001010011001010000000001000001000000010000110001000000000010101000000000000111100000000001000000100000110100001001100000000010000000000000000000011000000110000100100000100000100001000000000000000000001000010100000000000000000001100000001000100111010000001010010100010001111010100001000010101011000010100000000011100001000000110100001000000001000000000000000000100000110001001011001010000001000000010000000001001100001000001110000000000000001010000000010100001000011010000000001100000000000000000000000000000000001111000000010000000000011000000000100010100010010000000000000000000000001100110000001
// X3Y11, RegFile
`define Tile_X3Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000001100000000101100000000000000000000100000000000000000000000000000000000000010010110010100000000000000000000111000101110100001011001011100001100100010000000100101000000000000010000001001000000001011001100000000000000000000001000000000001010011101100011010100101001000000000010000001011101100000000000000000000100000001010000000000000010000000000000000011101100101011000011000000000000100000000000
// X4Y11, LUT4AB
`define Tile_X4Y11_Emulate_Bitstream 640'b0000001000000000000010100010000000011110101000000111001010000000000100100011010100000000001000000000000010000100000000000000010000011000100000110000000000000010000000010010000001000000000100000000000000000000010000000000001000000100000010000000000011000100000000111000101001000001110000100010010000100000000111101111011100001000001000000000100000010000000010000001000000100000100001000110000000000100001111010001010010010000110000001111000010000000000000000000000010000000000010001000010000101110000000001010100001000000100010000000000000000000000000011011010110010001001100000000000010000010000111110000010000000000010000010000001110010001
// X5Y11, LUT4AB
`define Tile_X5Y11_Emulate_Bitstream 640'b0000000000011010100010100000010000100110000001110000000010000000000000000011000000111110000000000000010000000000111100001010000000001000000000001010010000100011001010000000000000001100010000100001000110100000100100100010000100001000000010001000001000110001000000000000001100000000000101000000000000100000010101000000111000100000000000001010010000101000000000001000000000100001000001100111110100000001000000001001001110000000100001110010001100000000100000100000000100000000000000011010000001000100000000101000010001000000000010001100000011000000000000011101000111100010000000000000000100011000010000000000010000000000000000001001010010000000
// X6Y11, LUT4AB
`define Tile_X6Y11_Emulate_Bitstream 640'b0000000000000000101000001100000000000001110000000110000000001000000001000110100000010001000000000010000101111000000000100010000001100000000100010000000100100000000000000010000000100101111000000000010010000010010001001100001000000000000010001100110110010101001000000000000000000011000000000010000000000111000000000000110001011000000000100001100011100000100000000000000001000010000000001000000000011110011001100111101000010000000010010000100000000100000000000001010010100000000000000000000000100000001000000000000000000001000110010100000000010000000010010000010000001000001100000000001000000000000000001000000000000000100000000010000000000000
// X7Y11, DSP_top
`define Tile_X7Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000110000000000000000000000000000000000001010110000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000001100000000001011101110110000101100001101111010110000000000000000000000000000000000000000000011111101000000000000000011000000000000000000110000000010
// X8Y11, LUT4AB
`define Tile_X8Y11_Emulate_Bitstream 640'b0000000111100001011110000010000000000110000001110000000001111000001100000000110101100000000000100010000001000101011100000000000000100100000000001000100000010010000000000110000100000000110000000000000000000011110100010100000000000000000010000000001000100000000000011001100110001101000010010000000000010000000001101111010010011000011100000000000000010100010110001001000111001000100000000111000110010001010000010000100101001100010000010001110010100001100001100010010010000000001010010100101001000000001001010100010001000011000001010110000000110010000000001001100000001001001100000000000001100100110101000000000000000000100010000011010100010000
// X9Y11, LUT4AB
`define Tile_X9Y11_Emulate_Bitstream 640'b0000000000000110100011010010000000000010001000100110000001100000000000100001110001000000000000000001010000001001000000000000000000011000000000000100000100101011000000000000101001000000100011000000000000000000000000000000011000000010000100000000010010100000000000101100000000110001000000010011000001100001000000000000100100101000100110010000010011000000110001001001101011001011100000001000100001001111110100001100100000100000110011010001100100000000101001000000000001010000000010000000010000010001000001001001110001000000100000101000000000000000100000010000010001100001001000000000001000000011000000001010000000000000100001010010101010001000
// X10Y11, RAM_IO
`define Tile_X10Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000011000000000011111000000000000000000100001110100000000000000010000101000000000101010000011100000000100000000000000000010000000011110111110111110000000000000000100100101010101010101110101010110000001111100010100000001100111101010100100000111010011000001001
// X0Y12, W_IO
`define Tile_X0Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001110000000000000000000000
// X1Y12, LUT4AB
`define Tile_X1Y12_Emulate_Bitstream 640'b0000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000
// X2Y12, LUT4AB
`define Tile_X2Y12_Emulate_Bitstream 640'b0000000000000011000000100000000000011000110001000110000000000000000001000000110001100000000000000010000001011000000000000000000000000001000000000000000000100000000000000100100000100000100001000000000000100001010000001111000000000000000010010101000000000100001000010000110000100000000000000000000000011100100000001000001111000000011000000000001011010000110000001001000100001000100000001110000000000000001011011000010000011101010000000100101100010000000000100000000100010011010000000000010000000000011100001000100000000000000111101100000000000010000000011001010001000100001000000000000000000011011001000000000000000000100000001010000110001000
// X3Y12, RegFile
`define Tile_X3Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001100000100010001001000100000000101010000000000000000000000000000000110001001011110100000000000000000000011000000000110000000101011110001110100100010000001111110000000000010000000000110000100000100001000000000000000001000000110000000101011000000111001001011000100110111001111000100101101100001000011101010001001000000000011000010010010000000000010100000000000000000000000000000000000000111010
// X4Y12, LUT4AB
`define Tile_X4Y12_Emulate_Bitstream 640'b0000000000001110001001011000000000011110011000000011110000100000000001100101100010000111110010100000010000000010100100100111000000101001000000000110100000100100000000000000000100000000111100000000000010000100000110000000100101010000000000000000011010000110000000000001001101101000011001101000000000000000110000001111000100010000000011000010100100100101011010000000000000000000110000001001010100000000100001011000011000000000000000010100000100000001100000000000001111010000100010000100000001000100000000100011100000000010000100101100100010010000000000011111010001100000001100000000000010100101000000111000010000000000000000010101000100011000
// X5Y12, LUT4AB
`define Tile_X5Y12_Emulate_Bitstream 640'b0000000000001011101011110011110000000001111001000001001010000000000001101001000010100000000000000000000010010000101000000000000000000000000001110100000000010100001100000110000000001100101001100000000100101011100000000001101000000000000010000000000000001100001000000000001110000000000111110000000000000011000111000000010101100000001100001010000000101000011111000000000011101000000000001110100000011111001101001000101101000000000011000000000110001000000000100001100100010000000000000100000000110000001101010000100000000001010000011100100100000010000000010110010110001000001000000000001001011001011000000000000000000000100000111001001000001000
// X6Y12, LUT4AB
`define Tile_X6Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000011011000110001000000010000000000100001110000100000000000000000000000000000000100000000010000000000000000000000000000010001000000000110000001101100011000000000000000100101000000001111000000000000000010100000000000000000000000000000100100011001001111000000000000010001010100100000001110001000001001000000000011000000000111000001000111100000000000000000000000000000001000100000100001000000000000001000110100010001000000000001001000000000010000000000000001000110000010011000000100010000000100010000000111000010000101000100000001100000000000000000001100000000000000010000000000000000000000011000000000001000
// X7Y12, DSP_bot
`define Tile_X7Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000100000000000001001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000010000000000000000000000000000000000000111000000000000000000000000001000000011000001110000000000000000000000000111000000000000001000000000001001010000010000000000000000000000000000000000000000000000
// X8Y12, LUT4AB
`define Tile_X8Y12_Emulate_Bitstream 640'b0000001000000000100110001000100000000001100000000000010010101000000000000000000000000000000000000100000000000000000000010110000000000001100000100000100000000000010000001010010000000000001110000000010000010000000001111000000000000100000110100000100100000000000000001101100000100000100000000000010001000000000000010011010010000100010001001001110000000100010100000000001000001001101000000000000000011011010100000001001101011000000000010000010001000000000000100000100000000000000000000000010000000000000000110000000101000000000000011010001000000000000000010100000000111000000000001100001000000011000001110000000000000000111000101000101100101001
// X9Y12, LUT4AB
`define Tile_X9Y12_Emulate_Bitstream 640'b0000000000101110011000000000000000011111111001110000000000000000001101100111000000110000000000000001000000110000001000000110000001100000100000010000000000000000000000010000000000000000000000000000001100110000000010001000000000000000000000000000000011000000000000010000000000100001000100000000000000000001000000000100000010001100100000000000001000000000000000000001110001000001001000000000010000000100010100001000000000000001010010001000000110000000100010000000110000110000000101000000010000010000001000101000100100000000001000000000001000010000100000001101010000000001001100000101100000000000010001110000010000000000001100110101001010010010
// X10Y12, RAM_IO
`define Tile_X10Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110000000000000000100000000000000100000000000001000101111010000000000000000000000011000100010100010000000100000010000000000000000000000000000011101001110111110000000000000000100001101000010100111011011001010000100010000000000000101100111100100000111000100000000011000000
// X0Y13, W_IO
`define Tile_X0Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001110000000000000000000000
// X1Y13, LUT4AB
`define Tile_X1Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X2Y13, LUT4AB
`define Tile_X2Y13_Emulate_Bitstream 640'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000100000000000000000010000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000100000000000000000000010000001000000000010000000000000000000100011000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X3Y13, RegFile
`define Tile_X3Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000001010000000000000000000000000000000000000000000000000000001000010000100000000000000000000011000101011010100000101111100001000000000110100110100011000100000000101010000110011110000100010000000000000000000000000001100001000000001110101000000100000000000000000000001101001111100000000000000001000000000000000000000000111000000000111000000000000000000000000000000000000000000000000
// X4Y13, LUT4AB
`define Tile_X4Y13_Emulate_Bitstream 640'b0000000000000000111011000100100000000000000000000111000000000000000000000000100000010000000000000000000000001000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000010000100010000000000100000000000000000001000010000010000000000000100000000000011000000000
// X5Y13, LUT4AB
`define Tile_X5Y13_Emulate_Bitstream 640'b0000000000001000100001000000000000000000000000000000000001010000000000000000000000000010000000000000000000000000000000001000000001100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000001000000000000000000000000000000010000000000000000000001010000000001000000000000000000000000000000000000000010000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000011000011000000100000000000000000010000100000000000000010000010000000000000000000000001000000000000000000010000000000000000000110000000000000000
// X6Y13, LUT4AB
`define Tile_X6Y13_Emulate_Bitstream 640'b0000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000100000000010000000000000000000000000000011000001000000000000000000000000000000110000000000000000000000010010000000000000000000000000000000011010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000110010000000000000
// X7Y13, DSP_top
`define Tile_X7Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y13, LUT4AB
`define Tile_X8Y13_Emulate_Bitstream 640'b0000000000000000100001000011000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000100000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000010000000000001000000000000000000010000000000000010100000000000000000000000000000000010000000000000000000000000000000000100000000000000100000100110010000000000000000010000000000001000001000000000000000010000000000000000000000000000010000010000011010000000000000000000000000000001000000000000000000000000001000000000000000
// X9Y13, LUT4AB
`define Tile_X9Y13_Emulate_Bitstream 640'b0000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000100000100000000000000000000000000000000000000000100000100001000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000001000000000000001000000010000000000010000000000000000000010000001000010000
// X10Y13, RAM_IO
`define Tile_X10Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100010011000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000001000000000000000
// X0Y14, W_IO
`define Tile_X0Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001110000000000000000000000
// X1Y14, LUT4AB
`define Tile_X1Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X2Y14, LUT4AB
`define Tile_X2Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000
// X3Y14, RegFile
`define Tile_X3Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y14, LUT4AB
`define Tile_X4Y14_Emulate_Bitstream 640'b0000000000001011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000001000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000101000001000000000000000000000000000000001000000000
// X5Y14, LUT4AB
`define Tile_X5Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X6Y14, LUT4AB
`define Tile_X6Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X7Y14, DSP_bot
`define Tile_X7Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y14, LUT4AB
`define Tile_X8Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y14, LUT4AB
`define Tile_X9Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y14, RAM_IO
`define Tile_X10Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y15, W_IO
`define Tile_X0Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001110000000000000000000000
// X1Y15, LUT4AB
`define Tile_X1Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X2Y15, LUT4AB
`define Tile_X2Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X3Y15, RegFile
`define Tile_X3Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y15, LUT4AB
`define Tile_X4Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X5Y15, LUT4AB
`define Tile_X5Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X6Y15, LUT4AB
`define Tile_X6Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X7Y15, DSP_top
`define Tile_X7Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y15, LUT4AB
`define Tile_X8Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y15, LUT4AB
`define Tile_X9Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y15, RAM_IO
`define Tile_X10Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000
// X0Y16, W_IO
`define Tile_X0Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101111110000000000000000000000
// X1Y16, LUT4AB
`define Tile_X1Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000011111111000000000000000000000000001100111000000000000000000000000000000110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000
// X2Y16, LUT4AB
`define Tile_X2Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X3Y16, RegFile
`define Tile_X3Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y16, LUT4AB
`define Tile_X4Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X5Y16, LUT4AB
`define Tile_X5Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X6Y16, LUT4AB
`define Tile_X6Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X7Y16, DSP_bot
`define Tile_X7Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y16, LUT4AB
`define Tile_X8Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y16, LUT4AB
`define Tile_X9Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y16, RAM_IO
`define Tile_X10Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
