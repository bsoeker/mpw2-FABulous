// X0Y1, W_IO
`define Tile_X0Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y1, LUT4AB
`define Tile_X1Y1_Emulate_Bitstream 640'b0000000000000000010000110000000000000001010001110000000000000000000000110000010000000100000000100000010100000000000000000011000000000000000100010100100000010010001100000001000000001100001010000001100000000000010000001000111001011000000000000000000001001011001000000000000001000000000011001000000000000101000100001100000111111000000010001000000000001000011001000000000000100001100000100111110000000101100001001000000010000000000000100000000000000001100000000000000110010000000000001000000001000000010000000011000000000001000111000100000000000000000000001000001100100010000000000000000010000010000001110000000000000000000000000000001101000000
// X2Y1, LUT4AB
`define Tile_X2Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000100011001000000000000000000000000000100100000000000000000000000000000000000000001000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000110000000010000000000001000000000010000000000000000000110000000000000000101001000000000110000000000000000011000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000001000100100000000000000100010000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000
// X3Y1, RegFile
`define Tile_X3Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000011000000000000000100000000000000110000000010000000000000000000100000000000001110000000000000000000000000000000000000000000000000000
// X4Y1, LUT4AB
`define Tile_X4Y1_Emulate_Bitstream 640'b0000000000000000000100000000000000000001111000000111110000000000001000001111110001000010000000000100010000101001000000001000000000011000000110001101010100000000011010000010001100000000010000100001001000000001000010001000000101011010000000100001011001010010000000000000010011000110011001010000000000001010111100000011001010100000001000100000000000010000010001000000000000010000001001000000010000010000001100110000001010000000000011001100000101000001000000000000100000000000001000001000000001101100000000010001000100000011010110000100000010010000000000000000001001100000000100000000000010000000100010000000000000000000000000000000110100000000
// X5Y1, LUT4AB
`define Tile_X5Y1_Emulate_Bitstream 640'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000110000000000000000000000000100000100000000000000000001000000000000000100001000000011001001000010000100000000000000010000000000000010000000000000011001101010000001000000000000010000000000000000000000001000000000000000110000000010010000010001000000000000000000000011000000100000000000000100000001000000000001000000000000000010000010100000000000001000000000000000100000000000000000000000000000000100010000000000000000000000000000000000000000000000000001000000000000000000000
// X6Y1, LUT4AB
`define Tile_X6Y1_Emulate_Bitstream 640'b0000000000000000001000000010100000011001100000000000000000000000000001100011000000000000000000000000000000000000010100000000000000000000000000001110000000000010000000000000001000100000100000000000000000000000010000000000001000000000000000000100000000000000000000000000001101011000000001000000000000001101010000001100000000000000000000111000000000011000000000100000000000001110100001000000000000000000010000000000000000101000000011000000001000000000000000000000000000000000000000000000000000000010000010000000000000000000100000000000000000000000000000000000001000100100000000000000001000000000000111100000000000000000000000000000000000000000
// X7Y1, DSP_top
`define Tile_X7Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y1, LUT4AB
`define Tile_X8Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y1, LUT4AB
`define Tile_X9Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y1, RAM_IO
`define Tile_X10Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y2, W_IO
`define Tile_X0Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000110000000000000000000000000000000000000000000000000000000000000000
// X1Y2, LUT4AB
`define Tile_X1Y2_Emulate_Bitstream 640'b0000000000000000000000100000110000000000110001000000000000000000001001011000000010000000000000100000010001000000000000001001000001000000000100010110010000010000011000000010000000000001010010001000000100000000010100001001011011010001000010000100000011001011001000010000000001000001000011000000000010000001001000010000001011110000000010111000010000010000010001000000000001010010000001000111110000000000100000110000001000000000000000100011000100000000110000000000000010110000000000000000000001000100001100000011010000000000100001100000100000000000000000011001101000000011000000000000000000000000011101110010000000000000000000000000001001001010
// X2Y2, LUT4AB
`define Tile_X2Y2_Emulate_Bitstream 640'b0000000000000000111000101000100000000000000000000000001000010000000001100011100100000100000000100000000000000110100000100000000000001000100000001011110001010000000010010110001111000000101010100001111001000010110100101000101100001001001010110001110000000100001000000001101110001000000001001000000010010110010001011111000011000001001100100000010000010000011001000101000010100010001001100000000000010000001001001000100000010000110000110110000010000000101010100001000100110000100000000000010000011111100001001011000101000010100111000100000000010010000000010001001010000010000100000000000000000100100010010010010000000000000000000000000001100000
// X3Y2, RegFile
`define Tile_X3Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000110000000000000000000000001010000000000000010000010000000000011100100100000000000000000000000000011010001001110000000001110101000000000011010011001111000010101001000100000000001011000011010000000000000000000000000000000000000011001100000000000000001011101000001001001001010000000000001010000010101000011100000001000000001010000000110111000000000000000011000000001100000000000000000000
// X4Y2, LUT4AB
`define Tile_X4Y2_Emulate_Bitstream 640'b0000000000000001101000100010110000001110111001110001111000010000000001100100100001111100111110000000010000001010101100101010010000000001100000110110100000010000010000000001011000000001101010000000100000000111000000000100101000000010000010000000100000111001001001001000100101001010100100001010000000001101010100110000000111010000000000000000001100000100011111000000000001100110100001000000000000010111010000000010000001000000000011110000100000000100000100000001010000100000000000000000010001000010111100100010000001000011000000000000001000000000000000000010000000011000010000000000001111001000000001000001010000000000100100011000000000000000
// X5Y2, LUT4AB
`define Tile_X5Y2_Emulate_Bitstream 640'b0000000000000010010000100100000000000010001000000000010011010000001100100001100011100100000110100010000001000001000000000000010001000000000011101101010000010010010010000100010010000000100000000000010010001101000100000010000000000100000010100000000000110000000000000001101001000000000100000011000000001000011000001100000100000000000110100000001011001000000100000000000010010000100000100111000000010101101100000000000011000000000010001010100010000000100000100000000000100000000100011000010000001000010000000000010100000000000000001101000000000010000000011100001101001000000100000000001110000100000001100000000000000000000000000001001001100000
// X6Y2, LUT4AB
`define Tile_X6Y2_Emulate_Bitstream 640'b0000000000000000000000000001010000000000000000000000101000000000000000000000000000000000101000000000000001000001000001100000000000100000000110001001100000000000000000000000100000101000000000000000000100100000000000000100001100000100000000010000000010100000000000001000011000001000000010100010000000000010000010000000100000000000000100000000000000010000000011001000000000001010000000000000000100000000001000100000000000000000000000000000100000000000000000000000000001000000000000000100000000001010100000001010000000000001000100000000000000010000100000000110101000000000000100000000011000000100000111000000100000000000000000000001000000000000
// X7Y2, DSP_bot
`define Tile_X7Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000
// X8Y2, LUT4AB
`define Tile_X8Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y2, LUT4AB
`define Tile_X9Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y2, RAM_IO
`define Tile_X10Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y3, W_IO
`define Tile_X0Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y3, LUT4AB
`define Tile_X1Y3_Emulate_Bitstream 640'b0000000000000010010000000000000000010101010000000000000001111000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000100000000000000100000100000000010000000000000000000000000000000001000000000000010010000000000010000100000000010101100010000000010001110010000010001000000010000000010100000000000000100000000000001000000000000000000000000000000011000001000000000000000000011001110000000001010000000100000100000000000000000000000101000000000000001000000000001001010100110000000000010000000000000111100111100010000000000000001110000111000100000000000000000000000001001000000000000
// X2Y3, LUT4AB
`define Tile_X2Y3_Emulate_Bitstream 640'b0000000000000001001100010000000000000010001000010000000001110000000000111101000010110011000110000000100010001010101000011110000000001000000001110010010110000100000010010100000000000000001000000000000100100001000100000000001000000110000000011000100000101000000000000000110001000000010010100010001100000010001100001101101000011000000010000010011100100000100000000000001000110000100000001110010100010001101010110000101110000000000000110110100100000000000000000001011000100000001000001000000001001010000100000011010001000001000110000001000000010000000000010000100000000000000100000000000010011000011000011010000000000000000000000000110011100000
// X3Y3, RegFile
`define Tile_X3Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100010000010000000000000010000000111110000000000010000010000000000000011100000100000000000000000000000000011000100101001001100001111110001100010000000011001001110010101100110000000000010110000011010000000000010100010001000000000000000010010001100101011000111001001010000000001010111101101101001001001000000100000011110010000000000011010100000111001000000000000011000000000000000000000000000011
// X4Y3, LUT4AB
`define Tile_X4Y3_Emulate_Bitstream 640'b0000000000000110111000010000000000000001111000000000001010011000000000110101100001100001010010000001110110000000010100000011000000100001100000110001110011000011000010000100110010101001001110001000100010101001000100100101000010000100000010000001110000010000000000000000100000000001000100010000000000010001000000100011000000001000001101000000001000000100000111000000000001000010000000000001000100011111010010000000100101000000000011101000001000000000100000000000010000110000001000010000000001000100010010010000100100000001000010101101100000000000000000010010001101100000001000000000001000000100111001000010000000000000000000010110000100010000
// X5Y3, LUT4AB
`define Tile_X5Y3_Emulate_Bitstream 640'b0000000000000000100000000000100000000011101000000111001010011000000000110001000011110010000000000000000000010011111100011110000001000100100000110110000000001000010100000000001000000000100110100001100000000000000101000010001110001000000000000001100001000000000000000001100001100000000001000000000000000000001100010011001000001000001001100000001011100000000000000000000011010010100000000001000000001001001100000000100100100001000000100010101111010000011000100000000100100000010100000110000000101010011100010011100000000000011000010100000010000000000000010001000100001100001000000000001000000000001000000010000000000000000000101000000001010000
// X6Y3, LUT4AB
`define Tile_X6Y3_Emulate_Bitstream 640'b0000000000000000000011000010000000000000000001000110000000000000000000000000000000001100000100100000000001010110000001100000010001000000000110001000000101000100010010000000101010001100100100100000001100000000000110000001001000000100001000001101011010000000000000000000110010000010010010100010000000001001101110000011101000001000001000000000011100100001000000000000000000100000001100001000000000000000001000000000101000001000000000011000000000001001000000000000001000000000000100000000000000000100011010001100000100000000000000000010000000000000000000001101011000000100000100000000000000010011000010000000000000000000000000000010010011000010
// X7Y3, DSP_top
`define Tile_X7Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000100001100000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000001011000000000000000000000000000000000000
// X8Y3, LUT4AB
`define Tile_X8Y3_Emulate_Bitstream 640'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000
// X9Y3, LUT4AB
`define Tile_X9Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y3, RAM_IO
`define Tile_X10Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000
// X0Y4, W_IO
`define Tile_X0Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000
// X1Y4, LUT4AB
`define Tile_X1Y4_Emulate_Bitstream 640'b0000000000000000000000100000000000111111111001000110000000000000000000011000000110000001000000000000000100000110001000000010000000000000000110001100100100000000000000000000011001100000001010000000100000000000000100101100100100000000000000000000010000001000000010001000001000001000100010000000001100000010010001100100010100000000000000000000000000000000000011000000001000000000000000000110000000000100001000000000000000001000000010000000000000000000000000000000000000000000000000010000000000000000000010000011000000000001100101010100000000000000100000010100000100100100000000000000010100000000000011110000000000000000000000000000000010000000
// X2Y4, LUT4AB
`define Tile_X2Y4_Emulate_Bitstream 640'b0000000000000000010001011011100000100100111001111011110011101000000101110010000000010010000000100001110010000000111100000001000001010100100011110100010011111001000011010100100110000001100010100001000100001010000000000000010100001110000010000000010000101001110010000001100011100000111110100000101101010001010100000000101010000000010000001010001100010001110000001000000001000000010000001000010100010001010111000110010110001110000001010101101010000100101100000000000110010000000001000010010001100010000101101000010100000000100100010111100000000000000000010001011101101010000000000011101010000000100100010000100000000000000000000100110011110000
// X3Y4, RegFile
`define Tile_X3Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000100000000000000000001000100010000000000000000001000000000000001101000110110100000000000000000000111110101011100100000001110100100000000000001010100000110000000000010010110000000010110001000001000000000000000000100000001100000111011101010111000010110000001000101011101001010011100111100000000001111000000100000001000000000000010101100101000100000000000011000000000000000000000000001000
// X4Y4, LUT4AB
`define Tile_X4Y4_Emulate_Bitstream 640'b0000000000000000100000110000100000000001111000111001000000001000000000000000100000110001000000000000010000000000101000000010000000010000000000000010000000000000000100010001000010001000010000000001000111100101110001000000000000001000000000001100110000011000000000010001000001010111000110000000000000000001000101001000001100001000000000001011011100010001000110000010000001001000000000000111000000010110000000010000010101000000000011110010000100000000110100000000100000100000000000000000010000101000011100000000000100000001000000100001100010000010000000010000000001010001000000000000000101010010001000011010000000000000100000010000010001100000
// X5Y4, LUT4AB
`define Tile_X5Y4_Emulate_Bitstream 640'b0000000000000100110110110100000000100110011000110000000001111000001100000000000011100111001000000001010000000010010100011101010001000000100000000100000011000100010010000000001010001100000000000000100100000000000100001000000101010000000000000100001001000010000000000000000001000001000001100011000000000011001000111000000000000010000010011000011100100000000001010000000010010010100000101000000000000010110100100000001000001010000001110000000100000000010100000001000001000000100000010000010000001010100010000000100000000001000000000110000000000000000000011111000010000110000100000000001011101000010000010010100000000000000000000000101010000010
// X6Y4, LUT4AB
`define Tile_X6Y4_Emulate_Bitstream 640'b0000000000011000000000001100100000010110000000100100000000000000000100000010010001010000000000000010000000101110000000000000000000000001100000001000000100011010000100000000001001000000010101101001001000000110010000101001101111011000000000000100000000100000000000000000001110000000010010000000000000001101100010100011001010000000000000000000000000000000010010001000000001000010000000000111000000000100010010111000100010000100000001000000000100000000100100000001001000000001000000001000000000000110000000000000000000000000000100100000000000010000000010010000001010000011000100000000000000000000000000101010000000000000101000110100000000000010
// X7Y4, DSP_bot
`define Tile_X7Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000
// X8Y4, LUT4AB
`define Tile_X8Y4_Emulate_Bitstream 640'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000
// X9Y4, LUT4AB
`define Tile_X9Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y4, RAM_IO
`define Tile_X10Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000
// X0Y5, W_IO
`define Tile_X0Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000011000000000010000000000000000000000000000000000011000001100000000000000000000000
// X1Y5, LUT4AB
`define Tile_X1Y5_Emulate_Bitstream 640'b0000000000000000111000100000000000010001000000100000000000000000000100001010000101010010000000000110000110111101000100011100000000110001100100100000000100011000000000000000010100000000011100001000100100000010100000000000100010000000000100011000000001100000110000000001010111000000100000001000000000000000010010001111000010000000000000000000000100110000011000000000000000001010100001000001000000010000001010000000001000000000000000010101001000000001000000100001010000000000001000000000000001001100000011001001000000000010100000001000100000000010000000010101110000100000001100000000001010010000100100000010100000000000000000000000000011010010
// X2Y5, LUT4AB
`define Tile_X2Y5_Emulate_Bitstream 640'b0000000000000000100101000000100000011110000001000110000001011000000000000000010000000000101100000000000000000001000001110100010000001000100000001101000101000100000010000000001010101000010001100001000010000000000000100000000100001110000000000001001010000000000000010001000011100000000000111010000000000000111101000000011000001000000101000010011100100000101010000000000100010100100000001110000000000001011110110000001100010000000000000001000010000000000000000000000000100000000100010000010000001001101000000011000001000001100100000010000000010000000000011101000011011000001100000010000000010100010110010000000000000000000000100000010010001000
// X3Y5, RegFile
`define Tile_X3Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000010000000100010001000010010000000000000000000010001001011111000000000000000000000010010100101010111101001111001010000000000000000000000010000010000010000110000001100110000010000000000100000010000000000110000110000000001110000001000100000110110111010000011111001010100000000011101000100010000000010011000000000000000000011000000000000000000000000001100000000000000111000
// X4Y5, LUT4AB
`define Tile_X4Y5_Emulate_Bitstream 640'b0000000000000000000000001000000000000111111001010000001010011000000000010000000000100011000000000000010000010000001000000000000000000000000000010100010000000010010000110110001000000000011000000000000000001001110100001000000000000010000010101001000100000000000000011000000000001000000000000000000000000100000000010011000010010000001000100000001101100000010011000000000000000000000000000001000000010010000011000000011100000000000001011000000010000101000000100000000000000000001100000000000000101100000000011000000000000000000001000000000100000000100000000110001010101000000000000000000000101010110001111000010000000000000001001000000101000000
// X5Y5, LUT4AB
`define Tile_X5Y5_Emulate_Bitstream 640'b0000000000000010000110101110110000011001101001000110000011110000001100100000000000001111000110000011110100000000001000001000010000100101100000000000010000001011010010000000010011101000110100001000001100100111000001101110000011010100000010000000000101000000110000001000100000001001100001010010000000000000000101001100101000101000000000000000001111010001000011001000000000100000100000000110100000010001010000001000000000001100000000110010001010010000000000100000100000000000000000010000000001110000010001000000000000000000001010010110100010000000000000011010000010001011000000000000000011110000000000110000110000000000000000000000101001000010
// X6Y5, LUT4AB
`define Tile_X6Y5_Emulate_Bitstream 640'b0000000000010001011001110010000000001100110000000000000010001000000001100011000100000001000000100000000000000000000000000000000000001001100000000000000001001000000000000110000010001001100100100001000001000010000100000000000110001000001010100001000100000101001000000000100001001000011101010000000000010000010100001011000101000100000000011010000000100000000100000000000001100001100000000000010100010101000010100001011101000000000000001000000000000000000000000000001000110000000000000100000000000010000000000000100000000000000000010000000000000010000000000001000000000010001000000000000001001001100000100000000000000000000000010001000001000000
// X7Y5, DSP_top
`define Tile_X7Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000101000000000110000000000000000000000000000000000000000000000000000000000
// X8Y5, LUT4AB
`define Tile_X8Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y5, LUT4AB
`define Tile_X9Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y5, RAM_IO
`define Tile_X10Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y6, W_IO
`define Tile_X0Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110000000000000000000000000000000000000001101100010000000000000000000000000000000000000000000011100001110101000000000000000000
// X1Y6, LUT4AB
`define Tile_X1Y6_Emulate_Bitstream 640'b0000000000000000000000000000010000011110000000110001010000100000000000001000100001110011010010000000010001001001000000000000000000011000000111000000010100010100000000000000000000000000011000100000001110000000010100100000101001010110000000000101000110000001001000000001101100000000000001111000000000011110101001000000110101001000000100000000000100100100101010000000100110011001000000000001010000000011000110011000011000000000000000000001100100000000100000000001001000100000000000000000000000011000010100001001000000000001001100001100001000010000000100001001000100100010000000000100001100000100010000100000000000000000000000000010001000000000
// X2Y6, LUT4AB
`define Tile_X2Y6_Emulate_Bitstream 640'b0000000000000000000001000000010000010101010001010011111010000000000000000000100001000001000110000000010000000001000100000010010000000001000010000100100000010010001001000100110011000000001010000000100000000010100100001000101000000000000000101001010010000000000001010101000110000010100010001000001100011100010001010010010010101001000000001000010100000000011011010100100000000011100000000110111000010110010001000000100000010000000010000000000000000000001110100001000010000000000000000000010001010000011000000010000101000000000001000010000000000000000000001001010000011000000000000011000010110001011101000000100000000000000000000011000000000010
// X3Y6, RegFile
`define Tile_X3Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101001000000001000000000000000000000010000000000000000000000001000000000010000100111010101011110000010000000011110011100111000000101101110100001000000000000000001000000000000110000001100000000000011101111000000011100000011100000000000001010000010000000000000100110000000000010011000100000011011010000011001001000100000010001011011101101000000000111111100111011000011001100000000000000000000110000
// X4Y6, LUT4AB
`define Tile_X4Y6_Emulate_Bitstream 640'b0000000001100000111111000000000000100010001001111011001010101000000000100001000000011100001010100101010000000000011101100000000000010001100000001010110011000011010000000100101010001100000000100001000000000001100100001000001100001100000010001000010001110000000000010000001100010100000000000001000000000000000110000000000100101000000000001000000010101001010000000010100000101111100000100110100000010001000000000000011010000011100001001000000001000000001000100000001000000000000010011010010000010010000100000000010001000010000010000100000000010000000000000000001110000000011000000000001000011011000001000000110000000000100010010001100000000001
// X5Y6, LUT4AB
`define Tile_X5Y6_Emulate_Bitstream 640'b0000000000010000000100000000000000001011111000000000000000000000001001101001000000000000000000000010000101010000000000000000000000000000000100000000000000000100000001000000000000000000001010000000000000000000000000110001001000000000000000000000000010000001001000001000000000000001000000100000000000000000000100000000110101000000000000000010000000001000100000001000000001100000000000001000000000001101010000000000100000000000000000010000100010000000000000100000110000000000000000000000000011100000000001001010100000001000001000000010000010000000000000010010000111001000001000000000000000000001110100000000000000000000000000000000100000001000
// X6Y6, LUT4AB
`define Tile_X6Y6_Emulate_Bitstream 640'b0000000000000010011001100000000000011111100001110011011010111000000000000000100000101100011010000000010000010000101000001000010001001000000000010010000001100000000100000110000010000000110000100001001100000101000000000000100101011011000010100000010000010100001000001001101100000010010000000000000010000010001000000000111101010010001011000010001000000100100011001000000000010000000010001010011000010001110101101000000010000100000001110000100000001100000000000001010100110011001001001000000001111010010001101000010000000000000100000000101010000010000000000101000101100010000000000000000100000000110000000000000000000000000000011110000101010010
// X7Y6, DSP_bot
`define Tile_X7Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000110000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001001000000000000110000000000000000000000000000110000000000
// X8Y6, LUT4AB
`define Tile_X8Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000001000000000000000000000000000000001000000000000000000000000000111000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000001001000000000
// X9Y6, LUT4AB
`define Tile_X9Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000
// X10Y6, RAM_IO
`define Tile_X10Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000
// X0Y7, W_IO
`define Tile_X0Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100101111001000000000000000000
// X1Y7, LUT4AB
`define Tile_X1Y7_Emulate_Bitstream 640'b0000000000000010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000100000000000001000000000000000011000000010000000000000000000010000010010000010000000000000001000000010000000010010000000000000011000000011001000010000000000000000001000100000100110000000001001010000000000100000011100000000000000000100000000000000000000100001000000000000001000010001000010000000000000000000000001010000000000000000000000000000010011110000000000000000000000001000000001100001000000000000000000100000000110001000001000
// X2Y7, LUT4AB
`define Tile_X2Y7_Emulate_Bitstream 640'b0000000000000000011110100000100000000001111000100000101000000000000000001000100001001000101000000000010111001000000000000000000001000000000100000100110000001000010101000010001001000000011000000000000000101001000101100100100000000100000010000000000011100000000000000001100101001000000101001010000000000001001101001100111000000000001000100000001111000000001001000000001111010010100000000000000100010000001010000100001000000000110001000000000110001000011000100001110011000000000000010010000001001010000001100000000100000000010100000011000010010000100000000001011011000000001100000000010000000000110000111000000000000000000000001001101010001000
// X3Y7, RegFile
`define Tile_X3Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000001000000000111100000000010000000000000000000000000010100010001000000011000000000000011101011110001000000000000000000000111000000000110000110001101100010100010110110010100100000000100000110000001100100010101100010000000000000000000000000000001100001000000001110111101000101110001000000000011100000100000000011101010001101000011010110000101100001101010101110110000000000000111111000000000011000000000011000011
// X4Y7, LUT4AB
`define Tile_X4Y7_Emulate_Bitstream 640'b0000000000010110001001100000000000001010101000000000001010011000001100000000000000000011000110000110010100000000000000001000010000101000000000000100000010000111010000000111001010000001000001001000000000000111000000000011000010000010000010110000000010010100110000001001101111000000000001111011000000000101001000000000110000100010001010111000000011001000001000000000000001110101000000101111100001010110100011010001000010000110000001111001011010000000110000000101010101000000000000001001000000101101101100001011100010000000010111100000000000000000100000001011111101000101001000000000001010111001000010010000000000000000000001010010001001011000
// X5Y7, LUT4AB
`define Tile_X5Y7_Emulate_Bitstream 640'b0000000000001000110001100000100000000000000001111011110011111000000101100101000000010001000000100010010000000000001100000000000000000001100000000100000001010010000100000010000010001001001001001001100010001001000000001001101010001010000010000000010001100000000010000001110000010000100000001000100000000000010100110000100100001010001000001001101111101100001100000000000101000001000000000001001010011001010000000000001101010000000000101000001000000100100000000000000000010010000000000000000001001110000100000010010000000001000001001111100000000000000000000101010111110101001000000000000000011001001000010000000000000000100000001011000000001000
// X6Y7, LUT4AB
`define Tile_X6Y7_Emulate_Bitstream 640'b0000000000000100000000110010000000000000001001000110000000001000000000001000110001100101000000000000010000001000000000011000000000010000100000000101010000101000010100000100000010101001111110001001010100000000010100100111000000001100000010001100000000010010000000000000000001000001010000100000000000000100000100001100000110011000000010011111001000101100110000000000100000000110101000101111010010000000110000101000010010101001100000100001000000000001101000000000000000000000000000010000000000000000000010000000000100000101000100100000101000000000000000011101011010000110000100000000001010000001000001001000000000000000000000010000001000110000
// X7Y7, DSP_top
`define Tile_X7Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000010000000000000000000000000000000000000001110000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011000000000000000000110100000000000000000000000000000000
// X8Y7, LUT4AB
`define Tile_X8Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000110001000000000
// X9Y7, LUT4AB
`define Tile_X9Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y7, RAM_IO
`define Tile_X10Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010
// X0Y8, W_IO
`define Tile_X0Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000111100101110111000000000000000000
// X1Y8, LUT4AB
`define Tile_X1Y8_Emulate_Bitstream 640'b0000000000000000100101110000010000000000000000000000010011010000000000001000000110000100010100000001000010000000000000100000010000000000100111100010000001010000000000010110100000000000000011000000100000110110110000101010000000000100000000010001100000010100001000000000010000000000100100011001000000011100000000000011100001010001000100000000000000001000001000000100100000000000000000100110000100001001000100001000011100101000100000100000101110000000000000000000101001000000001100001100010000000110010101110011000000000010000100000100000000010010000000011010001000000110010000000000000100000101011001000010000000000000000000011000101010000010
// X2Y8, LUT4AB
`define Tile_X2Y8_Emulate_Bitstream 640'b0000000111000000001001000100100000001011001001010000000000000000000000100101000000100111110000000001000000000000001000000110000001101101100000010001010000000000000010110100100000000001011000001000010000100100010110101001001010000000000000100101100101001101111000010000001000001000000000000000000001011111100001001100011101000000000000001001100000000100000010000000000001000000110000000111000001001010000011001000010101000001000100110101000000010100100000000000101010010000000000010000010001010010001000010000100101000000110100000110000100110000100000001000101100100000001000000000001000000011101101111010010000000000000000001000000000111000
// X3Y8, RegFile
`define Tile_X3Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001010000011000000000000000000000001100000000100000000000000000000000110000000100010100000000000000000000111000000011110001000001110100011111110010001110100011110000000000000000001000010111000011000111000000000000000000000000000000001000100000001000000000000010000001100010001000100011100100001010011100000101010000001111110101100110010101111010010100000110000011000000000000000000000000000011
// X4Y8, LUT4AB
`define Tile_X4Y8_Emulate_Bitstream 640'b0000000000001011100101000101000000000110011001111011010011111000000100000000110000000011010110000000000000000000100000001000010000000000000000000010000001000010000100000001000011001000000100000001000000000000010000010000010100001100000000000100010111100010000000010000001100000000100000110000000000001100000100011011000000001000000000011000000001000000010000001000000001100000001000000110000100001100001011010000100000100100000000100101011000000000010000111000100010000000000000010000000000101101100101010000010001000000101100010000010100010000000000011101101101100000000000000010010001010000010100010010000000000000000000001001100000000000
// X5Y8, LUT4AB
`define Tile_X5Y8_Emulate_Bitstream 640'b0000000000000010000000101101010000001001100000100000000000001000001100001000000000010001000000000000010010010000000000000000000001001001000010000000000000000000010000000000110000000001111000001000110110000000000001111001000011000110000010000000000100000110000000000001100000001001000001000010000000000000001001010000010000001000000101000010000000010000010010001000000010111000000000000000000000010000000010100000000100011001000001110000000100000000001000000000010001000000000000000000000000011000100001011000100000000001101001000100000100000000000010000000000000000001001100000000001000000100011011000000000000000000000000001000001001010000
// X6Y8, LUT4AB
`define Tile_X6Y8_Emulate_Bitstream 640'b0000000000000000011111000000100000000000000000000000010010110000000100000000000100000000010010000001000010000100000000000000010000000000100000101000000001001110000000000000000101001000000001100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000111010000000000000010000100000100000000000000000000000000000000001101000001000000000000110000000001110000000000000000010000100000000001100000000000000110000001000000000000000010000000000000100000000000000000000010110010000000000000010000000010000010100000000000000010000100000100000100000000000000000000001001100101000000000000000000000000100100000000000
// X7Y8, DSP_bot
`define Tile_X7Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000001110111000000110000000011000000000000000000000000000000
// X8Y8, LUT4AB
`define Tile_X8Y8_Emulate_Bitstream 640'b0000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000011001000100000000
// X9Y8, LUT4AB
`define Tile_X9Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000
// X10Y8, RAM_IO
`define Tile_X10Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011111000000000000000000000000000001111010001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000011000010000000000110000000010
// X0Y9, W_IO
`define Tile_X0Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111110110000000000000000000
// X1Y9, LUT4AB
`define Tile_X1Y9_Emulate_Bitstream 640'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100001000000000000000000000000000000100001000000000000000000010001000000000000000000000000000000000000000000000000001000000000101000000000000000000000000000000000000100000000000000000110000000010000000000001000010100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000010000100000000000000000000000000001010000000100011000000000000000000000000000000000001000
// X2Y9, LUT4AB
`define Tile_X2Y9_Emulate_Bitstream 640'b0000000000000000000001111000000000001010101001110111000000000000000000000000110011100000000110000001000000000010100000011000010000110000000000000010000000001011001000000010000010000000001100001000001100000110010010011000000011010000000010100101100000000000000000010000001001000000000001010000000000010011100001010000000010110000000010011000011110010000010010000001000101000001000000000111110000010100100000101000000000000000010010101000000010000000000000100000000000000000000000010000010000001000011001000011100001000000000001000100000000000000000000001011110000000010001000000000000000000001010100001010000000000000000000000000001101000000
// X3Y9, RegFile
`define Tile_X3Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000111000000001000101011000000000000000000000000000000010110111000000000000000111000111001100001100010010111111000001100110110000000100000000000000000000000000000110000001011100000000000000010000000000010001100110101100000000111010110011010000001100110001000110110000011111110011100000111001000001011011100000000011000000100101000000000000010110000000000000000000000001000
// X4Y9, LUT4AB
`define Tile_X4Y9_Emulate_Bitstream 640'b0000000000000010110100010000010000000110111000000000101001000000000001100011000001001111000000000000010000001000011100001010010001100000000000001010010000110000010100110110000000101001110000000000000000100011010100100110000000000000000010000100010000110000000000000000101100000001000000000010000000010111011001001111110000000100001000011010010100100001100010000000000101010001000000101111000000010110000001000110101100010000110000100000000100001000010000100001111000000000100000000000000001101011100000000000000000000000000100010110100110010000000000001100000110000001000100000000001000000000100010010000000000000000000000010001101100010000
// X5Y9, LUT4AB
`define Tile_X5Y9_Emulate_Bitstream 640'b0000000000000000110010010000000000000000000001110011000010001000000000000000110001100000000000000000010000000000100001100000000001101100000000000110010000010010000100000000000100100000000000000001110000000000110010000100000000001000000000001100010000100000000000000000001000101110000011000000000000000010000000100000110000001000000100000000000010010000000001100010000000000010000000000000000000000100000000000000000000000000001010000000000001000100000100000000000000000000000000010000100001100000011110001000110000000010000000000000000000000000000000010000000010010100001000000000001001101100010000000000000000000000000000101001010010000001
// X6Y9, LUT4AB
`define Tile_X6Y9_Emulate_Bitstream 640'b0000000000001000010110000000000000000001111000000000011010111000000000000000000000000001010010000000010000000000000000010110010000000100000000000100000000010000010000000010000010001100011000000000100000000001000100000000000000000000000010000000100000110000000000000001000000000000101000000011000000000000000100010000111000000000000010000000000000000001000000000000000100001000000000000000010000010010100001100000010100000001001000000000000000000000011000000000000011000000000000000000000001000001100000000000000000000000000000000000000000010000000000010000101000000001000100000000000000000000100111000000000000000000000000010001100000011011
// X7Y9, DSP_top
`define Tile_X7Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000000000000000000101000000000000011010000000000000000000000000000000000000000000000000000
// X8Y9, LUT4AB
`define Tile_X8Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000001000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y9, LUT4AB
`define Tile_X9Y9_Emulate_Bitstream 640'b0000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000
// X10Y9, RAM_IO
`define Tile_X10Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000110001000000111000000000000000000000000101000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000010
// X0Y10, W_IO
`define Tile_X0Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y10, LUT4AB
`define Tile_X1Y10_Emulate_Bitstream 640'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000001000000000000000010000000000000000000000000110000100000000
// X2Y10, LUT4AB
`define Tile_X2Y10_Emulate_Bitstream 640'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000100000000000000000010000100000000000000000100000000000000000000000100000000000010000000000000000001000100000000110000000001000000001000000000000011000000000000000000000000000000000000000000011000000000000000000010000000010000000010000000001000000000000000000000100000000000000000000010000000000000000000000001000000000000001000000000000000000100000011000000000000000
// X3Y10, RegFile
`define Tile_X3Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000001000100000001000000101000000000101000001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y10, LUT4AB
`define Tile_X4Y10_Emulate_Bitstream 640'b0000000000000000000000100000000000000000101000110000000000000000000000000000100000100000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000001000000000001000000000000000000000001001010000000000000000010100000000000000010000000000000000000000000000000000000001000010000000000100000000000000000010000000000000000010000000000011000000000000000110000000000000000011000000000000000000000000000000000100000001000010000000000000000000000000000000000001000000011000011011000001000000000000001000100100010000000000010000000001100000100100000000001000000000100000010010000000000000000000000000000010000000
// X5Y10, LUT4AB
`define Tile_X5Y10_Emulate_Bitstream 640'b0000000000000001000000000010000000000000011000010000000000000000000000000000000000100001000000000000010000000000000000000000000000000000000000000010000000000000010000000010000000000000101000000000010000000000000100000000100000000000000010000000000000100010000000000000000100110000000001001000000001000000000000000000000100000000110000000011000000101000001000000000000001000000000000100000000000000000000001000000101010000001010000000000000000000000001000000000000010000000000000001000000000000000010000000000000000000000000000000000000000010010000000000010000000000000001000000000000000000000000110000010000000000000000000000000000000000000
// X6Y10, LUT4AB
`define Tile_X6Y10_Emulate_Bitstream 640'b0000000000000000100000000000000000000000000001010000000000001000000000000000000000000000000000000000010000000000000000000000000000001000100000100000000000000000000000000000000010000000000000000000001010100000000000000000010000000000000000000000000000000000000000000000000000000000000001100010000000000000000001000000010000000000000100000000100000010000000000001000000010001000001001000110000100000001000000000000100000000001010001000000100000000000001000000000000000000000000000000100010000000000010001001001000000000000000000000000010000010000000000000000100000010010000000000000001000000100000000000000000000000000000000000110000000000000
// X7Y10, DSP_bot
`define Tile_X7Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000001010000000000000000000000000000000000000000000000000000001100000000000000000000
// X8Y10, LUT4AB
`define Tile_X8Y10_Emulate_Bitstream 640'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000110000000000000000000000000000000010100000000000000000100000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000010010010000000000000000000000000000000000010001000000000000000000000000000000000000000000
// X9Y10, LUT4AB
`define Tile_X9Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000100100000000000010000000000000001000010000000000000100000000000000000000000000000000001000000000010000000000000000000000000100000000010000000000000000111000000000100000000000000000000000000000000100000000000000000000000000000000000000000
// X10Y10, RAM_IO
`define Tile_X10Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000001111000000000000000000001000000001010000000100000100000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000011100000000000
// X0Y11, W_IO
`define Tile_X0Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001100000000000000000000000
// X1Y11, LUT4AB
`define Tile_X1Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X2Y11, LUT4AB
`define Tile_X2Y11_Emulate_Bitstream 640'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000
// X3Y11, RegFile
`define Tile_X3Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000100000000000000000000000000110000000000000000000000000000000000000
// X4Y11, LUT4AB
`define Tile_X4Y11_Emulate_Bitstream 640'b0000000000000001000000001000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000110000000100000000000000000000000100000000000000000000000000100000000000100000001000000000010000100000000000000000000000000000010000000000100000000000010000000000000000000000000000000000000000000000000000001001100000000000100000100000000100000000000000100000000000010000000000000000010000000000000000010000000000000000000000011000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000
// X5Y11, LUT4AB
`define Tile_X5Y11_Emulate_Bitstream 640'b0000000000000101000111000000010000000000000000110000000000000000000000000000000001100000000000000000010000000000000000000000000000000000000000000100000000000010000000000000001001000000000000000000000100000000000000000000000000000000000110000000000010000000000000000001100000110001000000000000000000000000000010000000000000000000010001000000000000000000000001001000000010101000100000000110000000010000000100000000010100000000100001001000000110000000000001000000001000000000000000000001000000000000000001010000010010000000000000000010000100000010000000000000000000011001000000000011001000100000000000000000000000000000100000000110100000010000
// X6Y11, LUT4AB
`define Tile_X6Y11_Emulate_Bitstream 640'b0000000000000010000100000000100000000000000000110000000000000000000000000000000001100000000000000000000000000000000000000000000000000001100000100000000000000000000000100100010000100000000100000000000000000001000000000100011000000000000010000000000010000001001000000000000000100000000000000000010000000001000000000000000001000100000100000000000011000000000000101000000011000000000000000000000000010101001100101000001000000000000010000000000110000000000000000100000000010000001000000001000000000000000001000000000000000000000100000000010100000000000000001000000100000001100000000000000001110001000000000000000000000000100000000100101000011000
// X7Y11, DSP_top
`define Tile_X7Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010011000000100000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000001110101111000000000011110000000000000000000000000000000000000000000000000000000011010000000000000000000000000000000000000000
// X8Y11, LUT4AB
`define Tile_X8Y11_Emulate_Bitstream 640'b0000000000000100000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000101000000000000001000000000000010000000000000000000000010000000100000100000100000011000000000000100000000010000010000000000010000001100001001000100000000000000000000100000000000000000000000001000010000000000000100010000000011001000000000000000100000001000000000000000000000000000000000000000000010001000000000000000000000000000000000001000000000000000001100000000000000100001000
// X9Y11, LUT4AB
`define Tile_X9Y11_Emulate_Bitstream 640'b0000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000010000110000000000000000000000000000011100000000000000000000100000011100000000000000000000000000101111000000000000110000000000100000000000000011000000000000001001110001000010000000000110000000001100000011100000000000000101110010000000000000000000100010000001101101000000000000010010000001000011000000000000000000000000001000010000000000000000000000000010110111100000001000000001001000000011010100000000000000000000000000010000001000000001
// X10Y11, RAM_IO
`define Tile_X10Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100100111000000000000000000001000000000010000000000000000000000100001100000000000000000000100000010001000101000001000001000111110111011110010000000000000000000000000010101010011110001011110000001100000010001000000011111100000000100000001100010010001000
// X0Y12, W_IO
`define Tile_X0Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001110000000000000000000000
// X1Y12, LUT4AB
`define Tile_X1Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000
// X2Y12, LUT4AB
`define Tile_X2Y12_Emulate_Bitstream 640'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000
// X3Y12, RegFile
`define Tile_X3Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y12, LUT4AB
`define Tile_X4Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000010000
// X5Y12, LUT4AB
`define Tile_X5Y12_Emulate_Bitstream 640'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000001010000000
// X6Y12, LUT4AB
`define Tile_X6Y12_Emulate_Bitstream 640'b0000000000000101000001001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000010000000000100000000000000000000010000000000000010000000000000000000000000000001000000001000000000000000000000001000000100000000000000000000001000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001101000000000000000000000001000000010000000
// X7Y12, DSP_bot
`define Tile_X7Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001100000000000000000001000000001110000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000000000000000000001110000000001110000000000000000000001110000000000000011000000000000000001010000000000010000000000000000000000000000000010000000000000000000000000000000
// X8Y12, LUT4AB
`define Tile_X8Y12_Emulate_Bitstream 640'b0000000000000000011000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000100000000000000000000000000000001000000000000000000000000000000110001000000000001000000000000000001110010000000000100000010000000000011000000000000000000000000110000000101000000000000000000111110010001001100000000000000000000000010000000000000000001000000000000000000000010000000000000000000000000000000000000000100000000000000000000001000000000000001100000010010000000001000
// X9Y12, LUT4AB
`define Tile_X9Y12_Emulate_Bitstream 640'b0000000010011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000100100100000000000000000000000000100000010000000000100000000000000000000000000011001000000000001000000000001000010000000000100001000010101100000000000010010100011000000000000010000100000101000000001000000000000000000000000000010000000010000001000000000001001000000000000000100010000000000000000000000000000000011000
// X10Y12, RAM_IO
`define Tile_X10Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001010100000000000001000000000000000000000000000000001010001000011110000000000000000000100010100000000000000000000000000000100000100000000000000010001011111111101110000000000000000000010001010101000001010100110010000000000000000100000101111111100000000000000001010001011110000
// X0Y13, W_IO
`define Tile_X0Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001110000000000000000000000
// X1Y13, LUT4AB
`define Tile_X1Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X2Y13, LUT4AB
`define Tile_X2Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X3Y13, RegFile
`define Tile_X3Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y13, LUT4AB
`define Tile_X4Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X5Y13, LUT4AB
`define Tile_X5Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X6Y13, LUT4AB
`define Tile_X6Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X7Y13, DSP_top
`define Tile_X7Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000010100000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y13, LUT4AB
`define Tile_X8Y13_Emulate_Bitstream 640'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000
// X9Y13, LUT4AB
`define Tile_X9Y13_Emulate_Bitstream 640'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000010000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000001000000000010000000000000000000001000000000010000
// X10Y13, RAM_IO
`define Tile_X10Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000
// X0Y14, W_IO
`define Tile_X0Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001110000000000000000000000
// X1Y14, LUT4AB
`define Tile_X1Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X2Y14, LUT4AB
`define Tile_X2Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X3Y14, RegFile
`define Tile_X3Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y14, LUT4AB
`define Tile_X4Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X5Y14, LUT4AB
`define Tile_X5Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X6Y14, LUT4AB
`define Tile_X6Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X7Y14, DSP_bot
`define Tile_X7Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y14, LUT4AB
`define Tile_X8Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y14, LUT4AB
`define Tile_X9Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y14, RAM_IO
`define Tile_X10Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100
// X0Y15, W_IO
`define Tile_X0Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001110000000000000000000000
// X1Y15, LUT4AB
`define Tile_X1Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X2Y15, LUT4AB
`define Tile_X2Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X3Y15, RegFile
`define Tile_X3Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y15, LUT4AB
`define Tile_X4Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X5Y15, LUT4AB
`define Tile_X5Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X6Y15, LUT4AB
`define Tile_X6Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X7Y15, DSP_top
`define Tile_X7Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y15, LUT4AB
`define Tile_X8Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y15, LUT4AB
`define Tile_X9Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y15, RAM_IO
`define Tile_X10Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y16, W_IO
`define Tile_X0Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001110000000000000000000000
// X1Y16, LUT4AB
`define Tile_X1Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X2Y16, LUT4AB
`define Tile_X2Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X3Y16, RegFile
`define Tile_X3Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X4Y16, LUT4AB
`define Tile_X4Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X5Y16, LUT4AB
`define Tile_X5Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X6Y16, LUT4AB
`define Tile_X6Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X7Y16, DSP_bot
`define Tile_X7Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y16, LUT4AB
`define Tile_X8Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y16, LUT4AB
`define Tile_X9Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y16, RAM_IO
`define Tile_X10Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
